--******************************************************--
--        PONTIFICIA UNIVERSIDAD JAVERIANA              --
--                Disegno Digital                       --
--          Seccion de Tecnicas Digitales               --
-- 													              --
-- Titulo :    TestBenchModule                          --
-- Fecha  :  	D:XX M:XX Y:20XX                         --
--******************************************************--

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY TestProtocolRegisters IS
END TestProtocolRegisters;

ARCHITECTURE TestProtocolRegistersArch OF TestProtocolRegisters IS

--******************************************************--
-- Segnales a evaluar, las mismas definidas en el Work del bloque a evaluar
--******************************************************--

SIGNAL ControlSp        : STD_LOGIC_VECTOR( 1 DOWNTO 0) := "00";
SIGNAL ControlRegisters : STD_LOGIC_VECTOR(26 DOWNTO 0) := "000000000000000000000000000";
SIGNAL IrRegisters      : STD_LOGIC_VECTOR(31 DOWNTO 0) := x"00000000";
SIGNAL MemoryOut        : STD_LOGIC_VECTOR(31 DOWNTO 0) := x"00000000";
SIGNAL CsrRegisters     : STD_LOGIC_VECTOR(31 DOWNTO 0) := x"00000000";
SIGNAL AluRegisters     : STD_LOGIC_VECTOR(31 DOWNTO 0) := x"00000000";
SIGNAL PcRegisters      : STD_LOGIC_VECTOR(31 DOWNTO 0) := x"00000000";
SIGNAL Reset            : STD_LOGIC                     := '1';
SIGNAL Clk              : STD_LOGIC                     := '1';
SIGNAL RegistersCounter : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL MemoryIn         : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL RegistersMar     : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL RegistersCsr     : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL RegistersAlu     : STD_LOGIC_VECTOR(63 DOWNTO 0);

BEGIN

X58: ENTITY WORK.Registers 
PORT MAP	  (ControlSp        => ControlSp,
				ControlRegisters => ControlRegisters,
				IrRegisters      => IrRegisters,
				MemoryOut        => MemoryOut,
				CsrRegisters     => CsrRegisters,
				AluRegisters     => AluRegisters,
				PcRegisters      => PcRegisters,
				Reset            => Reset,
				Clk              => Clk,
				RegistersCounter => RegistersCounter,
				MemoryIn         => MemoryIn,
				RegistersMar     => RegistersMar,
				RegistersCsr     => RegistersCsr,
				RegistersAlu     => RegistersAlu
			  );

Clk   <= NOT Clk AFTER 10 ns;

Reset <= '0' AFTER 20 ns;

ControlSp <=   "00" AFTER 00020 ns,
					"00" AFTER 00040 ns,
					"00" AFTER 00060 ns,
					"00" AFTER 00080 ns,
					"00" AFTER 00100 ns,
					"00" AFTER 00120 ns,
					"00" AFTER 00140 ns,
					"00" AFTER 00160 ns,
					"00" AFTER 00180 ns,
					"00" AFTER 00200 ns,
					"00" AFTER 00220 ns,
					"00" AFTER 00240 ns,
					"00" AFTER 00260 ns,
					"00" AFTER 00280 ns,
					"00" AFTER 00300 ns,
					"00" AFTER 00320 ns,
					"00" AFTER 00340 ns,
					"00" AFTER 00360 ns,
					"00" AFTER 00380 ns,
					"00" AFTER 00400 ns,
					"00" AFTER 00420 ns,
					"00" AFTER 00440 ns,
					"00" AFTER 00460 ns,
					"00" AFTER 00480 ns,
					"00" AFTER 00500 ns,
					"00" AFTER 00520 ns,
					"00" AFTER 00540 ns,
					"00" AFTER 00560 ns,
					"00" AFTER 00580 ns,
					"00" AFTER 00600 ns,
					"00" AFTER 00620 ns,
					"00" AFTER 00640 ns,
					"00" AFTER 00660 ns,
					"00" AFTER 00680 ns,
					"00" AFTER 00700 ns,
					"00" AFTER 00720 ns,
					"00" AFTER 00740 ns,
					"00" AFTER 00760 ns,
					"00" AFTER 00780 ns,
					"00" AFTER 00800 ns,
					"00" AFTER 00820 ns,
					"00" AFTER 00840 ns,
					"00" AFTER 00860 ns,
					"00" AFTER 00880 ns,
					"00" AFTER 00900 ns,
					"00" AFTER 00920 ns,
					"00" AFTER 00940 ns,
					"00" AFTER 00960 ns,
					"00" AFTER 00980 ns,
					"00" AFTER 01000 ns,
					"00" AFTER 01020 ns,
					"00" AFTER 01040 ns,
					"00" AFTER 01060 ns,
					"00" AFTER 01080 ns,
					"00" AFTER 01100 ns,
					"00" AFTER 01120 ns,
					"00" AFTER 01140 ns,
					"00" AFTER 01160 ns,
					"00" AFTER 01180 ns,
					"00" AFTER 01200 ns,
					"00" AFTER 01220 ns,
					"00" AFTER 01240 ns,
					"00" AFTER 01260 ns,
					"00" AFTER 01280 ns,
					"00" AFTER 01300 ns,
					"00" AFTER 01320 ns,
					"00" AFTER 01340 ns,
					"00" AFTER 01360 ns,
					"00" AFTER 01380 ns,
					"00" AFTER 01400 ns,
					"00" AFTER 01420 ns,
					"00" AFTER 01440 ns,
					"00" AFTER 01460 ns,
					"00" AFTER 01480 ns,
					"00" AFTER 01500 ns,
					"00" AFTER 01520 ns,
					"00" AFTER 01540 ns,
					"00" AFTER 01560 ns,
					"00" AFTER 01580 ns,
					"00" AFTER 01600 ns,
					"00" AFTER 01620 ns,
					"00" AFTER 01640 ns,
					"00" AFTER 01660 ns,
					"00" AFTER 01680 ns,
					"00" AFTER 01700 ns,
					"00" AFTER 01720 ns,
					"00" AFTER 01740 ns,
					"00" AFTER 01760 ns,
					"00" AFTER 01780 ns,
					"00" AFTER 01800 ns,
					"00" AFTER 01820 ns,
					"00" AFTER 01840 ns,
					"00" AFTER 01860 ns,
					"00" AFTER 01880 ns,
					"00" AFTER 01900 ns,
					"00" AFTER 01920 ns,
					"00" AFTER 01940 ns,
					"00" AFTER 01960 ns,
					"00" AFTER 01980 ns,
					"00" AFTER 02000 ns,
					"00" AFTER 02020 ns,
					"00" AFTER 02040 ns,
					"00" AFTER 02060 ns,
					"00" AFTER 02080 ns,
					"00" AFTER 02100 ns,
					"00" AFTER 02120 ns,
					"00" AFTER 02140 ns,
					"00" AFTER 02160 ns,
					"00" AFTER 02180 ns,
					"00" AFTER 02200 ns,
					"00" AFTER 02220 ns,
					"00" AFTER 02240 ns,
					"00" AFTER 02260 ns,
					"00" AFTER 02280 ns,
					"00" AFTER 02300 ns,
					"00" AFTER 02320 ns,
					"00" AFTER 02340 ns,
					"00" AFTER 02360 ns,
					"00" AFTER 02380 ns,
					"00" AFTER 02400 ns,
					"00" AFTER 02420 ns,
					"00" AFTER 02440 ns,
					"00" AFTER 02460 ns,
					"00" AFTER 02480 ns,
					"00" AFTER 02500 ns,
					"00" AFTER 02520 ns,
					"00" AFTER 02540 ns,
					"00" AFTER 02560 ns,
					"00" AFTER 02580 ns,
					"00" AFTER 02600 ns,
					"00" AFTER 02620 ns,
					"00" AFTER 02640 ns,
					"00" AFTER 02660 ns,
					"00" AFTER 02680 ns,
					"00" AFTER 02700 ns,
					"00" AFTER 02720 ns,
					"00" AFTER 02740 ns,
					"00" AFTER 02760 ns,
					"00" AFTER 02780 ns,
					"00" AFTER 02800 ns,
					"00" AFTER 02820 ns,
					"00" AFTER 02840 ns,
					"00" AFTER 02860 ns,
					"00" AFTER 02880 ns,
					"00" AFTER 02900 ns,
					"00" AFTER 02920 ns,
					"00" AFTER 02940 ns,
					"00" AFTER 02960 ns,
					"00" AFTER 02980 ns,
					"00" AFTER 03000 ns,
					"00" AFTER 03020 ns,
					"00" AFTER 03040 ns,
					"00" AFTER 03060 ns,
					"00" AFTER 03080 ns,
					"00" AFTER 03100 ns,
					"00" AFTER 03120 ns,
					"00" AFTER 03140 ns,
					"00" AFTER 03160 ns,
					"00" AFTER 03180 ns,
					"00" AFTER 03200 ns,
					"00" AFTER 03220 ns,
					"00" AFTER 03240 ns,
					"00" AFTER 03260 ns,
					"00" AFTER 03280 ns,
					"00" AFTER 03300 ns,
					"00" AFTER 03320 ns,
					"00" AFTER 03340 ns,
					"00" AFTER 03360 ns,
					"00" AFTER 03380 ns,
					"00" AFTER 03400 ns,
					"00" AFTER 03420 ns,
					"00" AFTER 03440 ns,
					"00" AFTER 03460 ns,
					"00" AFTER 03480 ns,
					"00" AFTER 03500 ns,
					"00" AFTER 03520 ns,
					"00" AFTER 03540 ns,
					"00" AFTER 03560 ns,
					"00" AFTER 03580 ns,
					"00" AFTER 03600 ns,
					"00" AFTER 03620 ns,
					"00" AFTER 03640 ns,
					"00" AFTER 03660 ns,
					"00" AFTER 03680 ns,
					"00" AFTER 03700 ns,
					"00" AFTER 03720 ns,
					"00" AFTER 03740 ns,
					"00" AFTER 03760 ns,
					"00" AFTER 03780 ns,
					"00" AFTER 03800 ns,
					"00" AFTER 03820 ns,
					"00" AFTER 03840 ns,
					"00" AFTER 03860 ns,
					"00" AFTER 03880 ns,
					"00" AFTER 03900 ns,
					"00" AFTER 03920 ns,
					"00" AFTER 03940 ns,
					"00" AFTER 03960 ns,
					"00" AFTER 03980 ns,
					"00" AFTER 04000 ns,
					"00" AFTER 04020 ns,
					"00" AFTER 04040 ns,
					"00" AFTER 04060 ns,
					"00" AFTER 04080 ns,
					"00" AFTER 04100 ns,
					"00" AFTER 04120 ns,
					"00" AFTER 04140 ns,
					"00" AFTER 04160 ns,
					"00" AFTER 04180 ns,
					"00" AFTER 04200 ns,
					"00" AFTER 04220 ns,
					"00" AFTER 04240 ns,
					"00" AFTER 04260 ns,
					"00" AFTER 04280 ns,
					"00" AFTER 04300 ns,
					"00" AFTER 04320 ns,
					"00" AFTER 04340 ns,
					"00" AFTER 04360 ns,
					"00" AFTER 04380 ns,
					"00" AFTER 04400 ns,
					"00" AFTER 04420 ns,
					"00" AFTER 04440 ns,
					"00" AFTER 04460 ns,
					"00" AFTER 04480 ns,
					"00" AFTER 04500 ns,
					"00" AFTER 04520 ns,
					"00" AFTER 04540 ns,
					"00" AFTER 04560 ns,
					"00" AFTER 04580 ns,
					"00" AFTER 04600 ns,
					"00" AFTER 04620 ns,
					"00" AFTER 04640 ns,
					"00" AFTER 04660 ns,
					"00" AFTER 04680 ns,
					"00" AFTER 04700 ns,
					"00" AFTER 04720 ns,
					"00" AFTER 04740 ns,
					"00" AFTER 04760 ns,
					"00" AFTER 04780 ns,
					"00" AFTER 04800 ns,
					"00" AFTER 04820 ns,
					"00" AFTER 04840 ns,
					"00" AFTER 04860 ns,
					"00" AFTER 04880 ns,
					"00" AFTER 04900 ns,
					"00" AFTER 04920 ns,
					"00" AFTER 04940 ns,
					"00" AFTER 04960 ns,
					"00" AFTER 04980 ns,
					"00" AFTER 05000 ns,
					"00" AFTER 05020 ns,
					"00" AFTER 05040 ns,
					"00" AFTER 05060 ns,
					"00" AFTER 05080 ns,
					"00" AFTER 05100 ns,
					"00" AFTER 05120 ns,
					"00" AFTER 05140 ns,
					"00" AFTER 05160 ns,
					"00" AFTER 05180 ns,
					"00" AFTER 05200 ns,
					"00" AFTER 05220 ns,
					"00" AFTER 05240 ns,
					"00" AFTER 05260 ns,
					"00" AFTER 05280 ns,
					"00" AFTER 05300 ns,
					"00" AFTER 05320 ns,
					"00" AFTER 05340 ns,
					"00" AFTER 05360 ns,
					"00" AFTER 05380 ns,
					"00" AFTER 05400 ns,
					"00" AFTER 05420 ns,
					"00" AFTER 05440 ns,
					"00" AFTER 05460 ns,
					"00" AFTER 05480 ns,
					"00" AFTER 05500 ns,
					"00" AFTER 05520 ns,
					"00" AFTER 05540 ns,
					"00" AFTER 05560 ns,
					"00" AFTER 05580 ns,
					"00" AFTER 05600 ns,
					"00" AFTER 05620 ns,
					"00" AFTER 05640 ns,
					"00" AFTER 05660 ns,
					"00" AFTER 05680 ns,
					"00" AFTER 05700 ns,
					"00" AFTER 05720 ns,
					"00" AFTER 05740 ns,
					"00" AFTER 05760 ns,
					"00" AFTER 05780 ns,
					"00" AFTER 05800 ns,
					"00" AFTER 05820 ns,
					"00" AFTER 05840 ns,
					"00" AFTER 05860 ns,
					"00" AFTER 05880 ns,
					"00" AFTER 05900 ns,
					"00" AFTER 05920 ns,
					"00" AFTER 05940 ns,
					"00" AFTER 05960 ns,
					"00" AFTER 05980 ns,
					"00" AFTER 06000 ns,
					"00" AFTER 06020 ns,
					"00" AFTER 06040 ns,
					"00" AFTER 06060 ns,
					"00" AFTER 06080 ns,
					"00" AFTER 06100 ns,
					"00" AFTER 06120 ns,
					"00" AFTER 06140 ns,
					"00" AFTER 06160 ns,
					"00" AFTER 06180 ns,
					"00" AFTER 06200 ns,
					"00" AFTER 06220 ns,
					"00" AFTER 06240 ns,
					"00" AFTER 06260 ns,
					"00" AFTER 06280 ns,
					"00" AFTER 06300 ns,
					"00" AFTER 06320 ns,
					"00" AFTER 06340 ns,
					"00" AFTER 06360 ns,
					"00" AFTER 06380 ns,
					"00" AFTER 06400 ns,
					"00" AFTER 06420 ns,
					"00" AFTER 06440 ns,
					"00" AFTER 06460 ns,
					"00" AFTER 06480 ns,
					"00" AFTER 06500 ns,
					"00" AFTER 06520 ns,
					"00" AFTER 06540 ns,
					"00" AFTER 06560 ns,
					"00" AFTER 06580 ns,
					"00" AFTER 06600 ns,
					"00" AFTER 06620 ns,
					"00" AFTER 06640 ns,
					"00" AFTER 06660 ns,
					"00" AFTER 06680 ns,
					"00" AFTER 06700 ns,
					"00" AFTER 06720 ns,
					"00" AFTER 06740 ns,
					"00" AFTER 06760 ns,
					"00" AFTER 06780 ns,
					"00" AFTER 06800 ns,
					"00" AFTER 06820 ns,
					"00" AFTER 06840 ns,
					"00" AFTER 06860 ns,
					"00" AFTER 06880 ns,
					"00" AFTER 06900 ns,
					"00" AFTER 06920 ns,
					"00" AFTER 06940 ns,
					"00" AFTER 06960 ns,
					"00" AFTER 06980 ns,
					"00" AFTER 07000 ns,
					"00" AFTER 07020 ns,
					"00" AFTER 07040 ns,
					"00" AFTER 07060 ns,
					"00" AFTER 07080 ns,
					"00" AFTER 07100 ns,
					"00" AFTER 07120 ns,
					"00" AFTER 07140 ns,
					"00" AFTER 07160 ns,
					"00" AFTER 07180 ns,
					"00" AFTER 07200 ns,
					"00" AFTER 07220 ns,
					"00" AFTER 07240 ns,
					"00" AFTER 07260 ns,
					"00" AFTER 07280 ns,
					"00" AFTER 07300 ns,
					"00" AFTER 07320 ns,
					"00" AFTER 07340 ns,
					"00" AFTER 07360 ns,
					"00" AFTER 07380 ns,
					"00" AFTER 07400 ns,
					"00" AFTER 07420 ns,
					"00" AFTER 07440 ns,
					"00" AFTER 07460 ns,
					"00" AFTER 07480 ns,
					"00" AFTER 07500 ns,
					"00" AFTER 07520 ns,
					"00" AFTER 07540 ns,
					"00" AFTER 07560 ns,
					"00" AFTER 07580 ns,
					"00" AFTER 07600 ns,
					"00" AFTER 07620 ns,
					"00" AFTER 07640 ns,
					"00" AFTER 07660 ns,
					"00" AFTER 07680 ns,
					"00" AFTER 07700 ns,
					"00" AFTER 07720 ns,
					"00" AFTER 07740 ns,
					"00" AFTER 07760 ns,
					"00" AFTER 07780 ns,
					"00" AFTER 07800 ns,
					"00" AFTER 07820 ns,
					"00" AFTER 07840 ns,
					"00" AFTER 07860 ns,
					"00" AFTER 07880 ns,
					"00" AFTER 07900 ns,
					"00" AFTER 07920 ns,
					"00" AFTER 07940 ns,
					"00" AFTER 07960 ns,
					"00" AFTER 07980 ns,
					"00" AFTER 08000 ns,
					"00" AFTER 08020 ns,
					"00" AFTER 08040 ns,
					"00" AFTER 08060 ns,
					"00" AFTER 08080 ns,
					"00" AFTER 08100 ns,
					"00" AFTER 08120 ns,
					"00" AFTER 08140 ns,
					"00" AFTER 08160 ns,
					"00" AFTER 08180 ns,
					"00" AFTER 08200 ns,
					"00" AFTER 08220 ns,
					"00" AFTER 08240 ns,
					"00" AFTER 08260 ns,
					"00" AFTER 08280 ns,
					"00" AFTER 08300 ns,
					"00" AFTER 08320 ns,
					"00" AFTER 08340 ns,
					"00" AFTER 08360 ns,
					"00" AFTER 08380 ns,
					"00" AFTER 08400 ns,
					"00" AFTER 08420 ns,
					"00" AFTER 08440 ns,
					"00" AFTER 08460 ns,
					"00" AFTER 08480 ns,
					"00" AFTER 08500 ns,
					"00" AFTER 08520 ns,
					"00" AFTER 08540 ns,
					"00" AFTER 08560 ns,
					"00" AFTER 08580 ns,
					"00" AFTER 08600 ns,
					"00" AFTER 08620 ns,
					"00" AFTER 08640 ns,
					"00" AFTER 08660 ns,
					"00" AFTER 08680 ns,
					"00" AFTER 08700 ns,
					"00" AFTER 08720 ns,
					"00" AFTER 08740 ns,
					"00" AFTER 08760 ns,
					"00" AFTER 08780 ns,
					"00" AFTER 08800 ns,
					"00" AFTER 08820 ns,
					"00" AFTER 08840 ns,
					"00" AFTER 08860 ns,
					"00" AFTER 08880 ns,
					"00" AFTER 08900 ns,
					"00" AFTER 08920 ns,
					"00" AFTER 08940 ns,
					"00" AFTER 08960 ns,
					"00" AFTER 08980 ns,
					"00" AFTER 09000 ns,
					"00" AFTER 09020 ns,
					"00" AFTER 09040 ns,
					"00" AFTER 09060 ns,
					"00" AFTER 09080 ns,
					"00" AFTER 09100 ns,
					"00" AFTER 09120 ns,
					"00" AFTER 09140 ns,
					"00" AFTER 09160 ns,
					"00" AFTER 09180 ns,
					"00" AFTER 09200 ns,
					"00" AFTER 09220 ns,
					"00" AFTER 09240 ns,
					"00" AFTER 09260 ns,
					"00" AFTER 09280 ns,
					"00" AFTER 09300 ns,
					"00" AFTER 09320 ns,
					"00" AFTER 09340 ns,
					"00" AFTER 09360 ns,
					"00" AFTER 09380 ns,
					"00" AFTER 09400 ns,
					"00" AFTER 09420 ns,
					"00" AFTER 09440 ns,
					"00" AFTER 09460 ns,
					"00" AFTER 09480 ns,
					"00" AFTER 09500 ns,
					"00" AFTER 09520 ns,
					"00" AFTER 09540 ns,
					"00" AFTER 09560 ns,
					"00" AFTER 09580 ns,
					"00" AFTER 09600 ns,
					"00" AFTER 09620 ns,
					"00" AFTER 09640 ns,
					"00" AFTER 09660 ns,
					"00" AFTER 09680 ns,
					"00" AFTER 09700 ns,
					"00" AFTER 09720 ns,
					"00" AFTER 09740 ns,
					"00" AFTER 09760 ns,
					"00" AFTER 09780 ns,
					"00" AFTER 09800 ns,
					"00" AFTER 09820 ns,
					"00" AFTER 09840 ns,
					"00" AFTER 09860 ns,
					"00" AFTER 09880 ns,
					"00" AFTER 09900 ns,
					"00" AFTER 09920 ns,
					"00" AFTER 09940 ns,
					"00" AFTER 09960 ns,
					"00" AFTER 09980 ns,
					"00" AFTER 10000 ns,
					"00" AFTER 10020 ns,
					"00" AFTER 10040 ns,
					"00" AFTER 10060 ns,
					"00" AFTER 10080 ns,
					"00" AFTER 10100 ns,
					"00" AFTER 10120 ns,
					"00" AFTER 10140 ns,
					"00" AFTER 10160 ns,
					"00" AFTER 10180 ns,
					"00" AFTER 10200 ns,
					"00" AFTER 10220 ns,
					"00" AFTER 10240 ns,
					"00" AFTER 10260 ns,
					"00" AFTER 10280 ns,
					"00" AFTER 10300 ns,
					"00" AFTER 10320 ns,
					"00" AFTER 10340 ns,
					"00" AFTER 10360 ns,
					"00" AFTER 10380 ns,
					"00" AFTER 10400 ns,
					"00" AFTER 10420 ns,
					"00" AFTER 10440 ns,
					"00" AFTER 10460 ns,
					"00" AFTER 10480 ns,
					"00" AFTER 10500 ns,
					"00" AFTER 10520 ns,
					"00" AFTER 10540 ns,
					"00" AFTER 10560 ns,
					"00" AFTER 10580 ns,
					"00" AFTER 10600 ns,
					"00" AFTER 10620 ns,
					"00" AFTER 10640 ns,
					"00" AFTER 10660 ns,
					"00" AFTER 10680 ns,
					"00" AFTER 10700 ns,
					"00" AFTER 10720 ns,
					"00" AFTER 10740 ns,
					"00" AFTER 10760 ns,
					"00" AFTER 10780 ns,
					"00" AFTER 10800 ns,
					"00" AFTER 10820 ns,
					"00" AFTER 10840 ns,
					"00" AFTER 10860 ns,
					"00" AFTER 10880 ns,
					"00" AFTER 10900 ns,
					"00" AFTER 10920 ns,
					"00" AFTER 10940 ns,
					"00" AFTER 10960 ns,
					"00" AFTER 10980 ns,
					"00" AFTER 11000 ns,
					"00" AFTER 11020 ns,
					"00" AFTER 11040 ns,
					"00" AFTER 11060 ns,
					"00" AFTER 11080 ns,
					"00" AFTER 11100 ns,
					"00" AFTER 11120 ns,
					"00" AFTER 11140 ns,
					"00" AFTER 11160 ns,
					"00" AFTER 11180 ns,
					"00" AFTER 11200 ns,
					"00" AFTER 11220 ns,
					"00" AFTER 11240 ns,
					"00" AFTER 11260 ns,
					"00" AFTER 11280 ns,
					"00" AFTER 11300 ns,
					"00" AFTER 11320 ns,
					"00" AFTER 11340 ns,
					"00" AFTER 11360 ns,
					"00" AFTER 11380 ns,
					"00" AFTER 11400 ns,
					"00" AFTER 11420 ns,
					"00" AFTER 11440 ns,
					"00" AFTER 11460 ns,
					"00" AFTER 11480 ns,
					"00" AFTER 11500 ns,
					"00" AFTER 11520 ns,
					"00" AFTER 11540 ns,
					"00" AFTER 11560 ns,
					"00" AFTER 11580 ns,
					"00" AFTER 11600 ns,
					"00" AFTER 11620 ns,
					"00" AFTER 11640 ns,
					"00" AFTER 11660 ns,
					"00" AFTER 11680 ns,
					"00" AFTER 11700 ns,
					"00" AFTER 11720 ns,
					"00" AFTER 11740 ns,
					"00" AFTER 11760 ns,
					"00" AFTER 11780 ns,
					"00" AFTER 11800 ns,
					"00" AFTER 11820 ns,
					"00" AFTER 11840 ns,
					"00" AFTER 11860 ns,
					"00" AFTER 11880 ns,
					"00" AFTER 11900 ns,
					"00" AFTER 11920 ns,
					"00" AFTER 11940 ns,
					"00" AFTER 11960 ns,
					"00" AFTER 11980 ns,
					"00" AFTER 12000 ns,
					"00" AFTER 12020 ns,
					"00" AFTER 12040 ns,
					"00" AFTER 12060 ns,
					"00" AFTER 12080 ns,
					"00" AFTER 12100 ns,
					"00" AFTER 12120 ns,
					"00" AFTER 12140 ns,
					"00" AFTER 12160 ns,
					"00" AFTER 12180 ns,
					"00" AFTER 12200 ns,
					"00" AFTER 12220 ns,
					"00" AFTER 12240 ns,
					"00" AFTER 12260 ns,
					"00" AFTER 12280 ns,
					"00" AFTER 12300 ns,
					"00" AFTER 12320 ns,
					"00" AFTER 12340 ns,
					"00" AFTER 12360 ns,
					"00" AFTER 12380 ns,
					"00" AFTER 12400 ns,
					"00" AFTER 12420 ns,
					"00" AFTER 12440 ns,
					"00" AFTER 12460 ns,
					"00" AFTER 12480 ns,
					"00" AFTER 12500 ns,
					"00" AFTER 12520 ns,
					"00" AFTER 12540 ns,
					"00" AFTER 12560 ns,
					"00" AFTER 12580 ns,
					"00" AFTER 12600 ns,
					"00" AFTER 12620 ns,
					"00" AFTER 12640 ns,
					"00" AFTER 12660 ns,
					"00" AFTER 12680 ns,
					"00" AFTER 12700 ns,
					"00" AFTER 12720 ns,
					"00" AFTER 12740 ns,
					"00" AFTER 12760 ns,
					"00" AFTER 12780 ns,
					"00" AFTER 12800 ns,
					"00" AFTER 12820 ns,
					"00" AFTER 12840 ns,
					"00" AFTER 12860 ns,
					"00" AFTER 12880 ns,
					"00" AFTER 12900 ns,
					"00" AFTER 12920 ns,
					"00" AFTER 12940 ns,
					"00" AFTER 12960 ns,
					"00" AFTER 12980 ns,
					"00" AFTER 13000 ns,
					"00" AFTER 13020 ns,
					"00" AFTER 13040 ns,
					"00" AFTER 13060 ns,
					"00" AFTER 13080 ns,
					"00" AFTER 13100 ns,
					"00" AFTER 13120 ns,
					"00" AFTER 13140 ns,
					"00" AFTER 13160 ns,
					"00" AFTER 13180 ns,
					"00" AFTER 13200 ns,
					"00" AFTER 13220 ns,
					"00" AFTER 13240 ns,
					"00" AFTER 13260 ns,
					"00" AFTER 13280 ns,
					"00" AFTER 13300 ns,
					"00" AFTER 13320 ns,
					"00" AFTER 13340 ns,
					"00" AFTER 13360 ns,
					"00" AFTER 13380 ns,
					"00" AFTER 13400 ns,
					"00" AFTER 13420 ns,
					"00" AFTER 13440 ns,
					"00" AFTER 13460 ns,
					"00" AFTER 13480 ns,
					"00" AFTER 13500 ns,
					"00" AFTER 13520 ns,
					"00" AFTER 13540 ns,
					"00" AFTER 13560 ns,
					"00" AFTER 13580 ns,
					"00" AFTER 13600 ns,
					"00" AFTER 13620 ns,
					"00" AFTER 13640 ns,
					"00" AFTER 13660 ns,
					"00" AFTER 13680 ns,
					"00" AFTER 13700 ns,
					"00" AFTER 13720 ns,
					"00" AFTER 13740 ns,
					"00" AFTER 13760 ns,
					"00" AFTER 13780 ns,
					"00" AFTER 13800 ns,
					"00" AFTER 13820 ns,
					"00" AFTER 13840 ns,
					"00" AFTER 13860 ns,
					"00" AFTER 13880 ns,
					"00" AFTER 13900 ns,
					"00" AFTER 13920 ns,
					"00" AFTER 13940 ns,
					"00" AFTER 13960 ns,
					"00" AFTER 13980 ns,
					"00" AFTER 14000 ns,
					"00" AFTER 14020 ns,
					"00" AFTER 14040 ns,
					"00" AFTER 14060 ns,
					"00" AFTER 14080 ns,
					"00" AFTER 14100 ns,
					"00" AFTER 14120 ns,
					"00" AFTER 14140 ns,
					"00" AFTER 14160 ns,
					"00" AFTER 14180 ns,
					"00" AFTER 14200 ns,
					"00" AFTER 14220 ns,
					"00" AFTER 14240 ns,
					"00" AFTER 14260 ns,
					"00" AFTER 14280 ns,
					"00" AFTER 14300 ns,
					"00" AFTER 14320 ns,
					"00" AFTER 14340 ns,
					"00" AFTER 14360 ns,
					"00" AFTER 14380 ns,
					"00" AFTER 14400 ns,
					"00" AFTER 14420 ns,
					"00" AFTER 14440 ns,
					"00" AFTER 14460 ns,
					"00" AFTER 14480 ns,
					"00" AFTER 14500 ns,
					"00" AFTER 14520 ns,
					"00" AFTER 14540 ns,
					"00" AFTER 14560 ns,
					"00" AFTER 14580 ns,
					"00" AFTER 14600 ns,
					"00" AFTER 14620 ns,
					"00" AFTER 14640 ns,
					"00" AFTER 14660 ns,
					"00" AFTER 14680 ns,
					"00" AFTER 14700 ns,
					"00" AFTER 14720 ns,
					"00" AFTER 14740 ns,
					"00" AFTER 14760 ns,
					"00" AFTER 14780 ns,
					"00" AFTER 14800 ns,
					"00" AFTER 14820 ns,
					"00" AFTER 14840 ns,
					"00" AFTER 14860 ns,
					"00" AFTER 14880 ns,
					"00" AFTER 14900 ns,
					"00" AFTER 14920 ns,
					"00" AFTER 14940 ns,
					"00" AFTER 14960 ns,
					"00" AFTER 14980 ns,
					"00" AFTER 15000 ns,
					"00" AFTER 15020 ns,
					"00" AFTER 15040 ns,
					"00" AFTER 15060 ns,
					"00" AFTER 15080 ns,
					"00" AFTER 15100 ns,
					"00" AFTER 15120 ns,
					"00" AFTER 15140 ns,
					"00" AFTER 15160 ns,
					"00" AFTER 15180 ns,
					"00" AFTER 15200 ns,
					"00" AFTER 15220 ns,
					"00" AFTER 15240 ns,
					"00" AFTER 15260 ns,
					"00" AFTER 15280 ns,
					"00" AFTER 15300 ns,
					"00" AFTER 15320 ns,
					"00" AFTER 15340 ns,
					"00" AFTER 15360 ns,
					"00" AFTER 15380 ns,
					"00" AFTER 15400 ns,
					"00" AFTER 15420 ns,
					"00" AFTER 15440 ns,
					"00" AFTER 15460 ns,
					"00" AFTER 15480 ns,
					"00" AFTER 15500 ns,
					"00" AFTER 15520 ns,
					"00" AFTER 15540 ns,
					"00" AFTER 15560 ns,
					"00" AFTER 15580 ns,
					"00" AFTER 15600 ns,
					"00" AFTER 15620 ns,
					"00" AFTER 15640 ns,
					"00" AFTER 15660 ns,
					"00" AFTER 15680 ns,
					"00" AFTER 15700 ns,
					"00" AFTER 15720 ns,
					"00" AFTER 15740 ns,
					"00" AFTER 15760 ns,
					"00" AFTER 15780 ns,
					"00" AFTER 15800 ns,
					"00" AFTER 15820 ns,
					"00" AFTER 15840 ns,
					"00" AFTER 15860 ns,
					"00" AFTER 15880 ns,
					"00" AFTER 15900 ns,
					"00" AFTER 15920 ns,
					"00" AFTER 15940 ns,
					"00" AFTER 15960 ns,
					"00" AFTER 15980 ns,
					"00" AFTER 16000 ns,
					"00" AFTER 16020 ns,
					"00" AFTER 16040 ns,
					"00" AFTER 16060 ns,
					"00" AFTER 16080 ns,
					"00" AFTER 16100 ns,
					"00" AFTER 16120 ns,
					"00" AFTER 16140 ns,
					"00" AFTER 16160 ns,
					"00" AFTER 16180 ns,
					"00" AFTER 16200 ns,
					"00" AFTER 16220 ns,
					"00" AFTER 16240 ns,
					"00" AFTER 16260 ns,
					"00" AFTER 16280 ns,
					"00" AFTER 16300 ns,
					"00" AFTER 16320 ns,
					"00" AFTER 16340 ns,
					"00" AFTER 16360 ns,
					"00" AFTER 16380 ns,
					"00" AFTER 16400 ns,
					"00" AFTER 16420 ns,
					"00" AFTER 16440 ns,
					"00" AFTER 16460 ns,
					"00" AFTER 16480 ns,
					"00" AFTER 16500 ns,
					"00" AFTER 16520 ns,
					"00" AFTER 16540 ns,
					"00" AFTER 16560 ns,
					"00" AFTER 16580 ns,
					"00" AFTER 16600 ns,
					"00" AFTER 16620 ns,
					"00" AFTER 16640 ns,
					"00" AFTER 16660 ns,
					"00" AFTER 16680 ns,
					"00" AFTER 16700 ns,
					"00" AFTER 16720 ns,
					"00" AFTER 16740 ns,
					"00" AFTER 16760 ns,
					"00" AFTER 16780 ns,
					"00" AFTER 16800 ns,
					"00" AFTER 16820 ns,
					"00" AFTER 16840 ns,
					"00" AFTER 16860 ns,
					"00" AFTER 16880 ns,
					"00" AFTER 16900 ns,
					"00" AFTER 16920 ns,
					"00" AFTER 16940 ns,
					"00" AFTER 16960 ns,
					"00" AFTER 16980 ns,
					"00" AFTER 17000 ns,
					"00" AFTER 17020 ns,
					"00" AFTER 17040 ns,
					"00" AFTER 17060 ns,
					"00" AFTER 17080 ns,
					"00" AFTER 17100 ns,
					"00" AFTER 17120 ns,
					"00" AFTER 17140 ns,
					"00" AFTER 17160 ns,
					"00" AFTER 17180 ns,
					"00" AFTER 17200 ns,
					"00" AFTER 17220 ns,
					"00" AFTER 17240 ns,
					"00" AFTER 17260 ns,
					"00" AFTER 17280 ns,
					"00" AFTER 17300 ns,
					"00" AFTER 17320 ns,
					"00" AFTER 17340 ns,
					"00" AFTER 17360 ns,
					"00" AFTER 17380 ns,
					"00" AFTER 17400 ns,
					"00" AFTER 17420 ns,
					"00" AFTER 17440 ns,
					"00" AFTER 17460 ns,
					"00" AFTER 17480 ns,
					"00" AFTER 17500 ns,
					"00" AFTER 17520 ns,
					"00" AFTER 17540 ns,
					"00" AFTER 17560 ns,
					"00" AFTER 17580 ns,
					"00" AFTER 17600 ns,
					"00" AFTER 17620 ns,
					"00" AFTER 17640 ns,
					"00" AFTER 17660 ns,
					"00" AFTER 17680 ns,
					"00" AFTER 17700 ns,
					"00" AFTER 17720 ns,
					"00" AFTER 17740 ns,
					"00" AFTER 17760 ns,
					"00" AFTER 17780 ns,
					"00" AFTER 17800 ns,
					"00" AFTER 17820 ns,
					"00" AFTER 17840 ns,
					"00" AFTER 17860 ns,
					"00" AFTER 17880 ns,
					"00" AFTER 17900 ns,
					"00" AFTER 17920 ns,
					"00" AFTER 17940 ns,
					"00" AFTER 17960 ns,
					"00" AFTER 17980 ns,
					"00" AFTER 18000 ns,
					"00" AFTER 18020 ns,
					"00" AFTER 18040 ns,
					"00" AFTER 18060 ns,
					"00" AFTER 18080 ns,
					"00" AFTER 18100 ns,
					"00" AFTER 18120 ns,
					"00" AFTER 18140 ns,
					"00" AFTER 18160 ns,
					"00" AFTER 18180 ns,
					"00" AFTER 18200 ns,
					"00" AFTER 18220 ns,
					"00" AFTER 18240 ns,
					"00" AFTER 18260 ns,
					"00" AFTER 18280 ns,
					"00" AFTER 18300 ns,
					"00" AFTER 18320 ns,
					"00" AFTER 18340 ns,
					"00" AFTER 18360 ns,
					"00" AFTER 18380 ns,
					"00" AFTER 18400 ns,
					"00" AFTER 18420 ns,
					"00" AFTER 18440 ns,
					"00" AFTER 18460 ns,
					"00" AFTER 18480 ns,
					"00" AFTER 18500 ns,
					"00" AFTER 18520 ns,
					"00" AFTER 18540 ns,
					"00" AFTER 18560 ns,
					"00" AFTER 18580 ns,
					"00" AFTER 18600 ns,
					"00" AFTER 18620 ns,
					"00" AFTER 18640 ns,
					"00" AFTER 18660 ns,
					"00" AFTER 18680 ns,
					"00" AFTER 18700 ns,
					"00" AFTER 18720 ns,
					"00" AFTER 18740 ns,
					"00" AFTER 18760 ns,
					"00" AFTER 18780 ns,
					"00" AFTER 18800 ns,
					"00" AFTER 18820 ns,
					"00" AFTER 18840 ns,
					"00" AFTER 18860 ns,
					"00" AFTER 18880 ns,
					"00" AFTER 18900 ns,
					"00" AFTER 18920 ns,
					"00" AFTER 18940 ns,
					"00" AFTER 18960 ns,
					"00" AFTER 18980 ns,
					"00" AFTER 19000 ns,
					"00" AFTER 19020 ns,
					"00" AFTER 19040 ns,
					"00" AFTER 19060 ns,
					"00" AFTER 19080 ns,
					"00" AFTER 19100 ns,
					"00" AFTER 19120 ns,
					"00" AFTER 19140 ns,
					"00" AFTER 19160 ns,
					"00" AFTER 19180 ns,
					"00" AFTER 19200 ns,
					"00" AFTER 19220 ns,
					"00" AFTER 19240 ns,
					"00" AFTER 19260 ns,
					"00" AFTER 19280 ns,
					"00" AFTER 19300 ns,
					"00" AFTER 19320 ns,
					"00" AFTER 19340 ns,
					"00" AFTER 19360 ns,
					"00" AFTER 19380 ns,
					"00" AFTER 19400 ns,
					"00" AFTER 19420 ns,
					"00" AFTER 19440 ns,
					"00" AFTER 19460 ns,
					"00" AFTER 19480 ns,
					"00" AFTER 19500 ns,
					"00" AFTER 19520 ns,
					"00" AFTER 19540 ns,
					"00" AFTER 19560 ns,
					"00" AFTER 19580 ns,
					"00" AFTER 19600 ns,
					"00" AFTER 19620 ns,
					"00" AFTER 19640 ns,
					"00" AFTER 19660 ns,
					"00" AFTER 19680 ns,
					"00" AFTER 19700 ns,
					"00" AFTER 19720 ns,
					"00" AFTER 19740 ns,
					"00" AFTER 19760 ns,
					"00" AFTER 19780 ns,
					"00" AFTER 19800 ns,
					"00" AFTER 19820 ns,
					"00" AFTER 19840 ns,
					"00" AFTER 19860 ns,
					"00" AFTER 19880 ns,
					"00" AFTER 19900 ns,
					"00" AFTER 19920 ns,
					"00" AFTER 19940 ns,
					"00" AFTER 19960 ns,
					"00" AFTER 19980 ns,
					"00" AFTER 20000 ns,
					"00" AFTER 20020 ns,
					"00" AFTER 20040 ns,
					"00" AFTER 20060 ns,
					"00" AFTER 20080 ns,
					"00" AFTER 20100 ns,
					"00" AFTER 20120 ns,
					"00" AFTER 20140 ns,
					"00" AFTER 20160 ns,
					"00" AFTER 20180 ns,
					"00" AFTER 20200 ns,
					"00" AFTER 20220 ns,
					"00" AFTER 20240 ns,
					"00" AFTER 20260 ns,
					"00" AFTER 20280 ns,
					"00" AFTER 20300 ns,
					"00" AFTER 20320 ns,
					"00" AFTER 20340 ns,
					"00" AFTER 20360 ns,
					"00" AFTER 20380 ns,
					"00" AFTER 20400 ns,
					"00" AFTER 20420 ns,
					"00" AFTER 20440 ns,
					"00" AFTER 20460 ns,
					"00" AFTER 20480 ns,
					"00" AFTER 20500 ns,
					"00" AFTER 20520 ns,
					"00" AFTER 20540 ns,
					"00" AFTER 20560 ns,
					"00" AFTER 20580 ns,
					"00" AFTER 20600 ns,
					"00" AFTER 20620 ns,
					"00" AFTER 20640 ns,
					"00" AFTER 20660 ns,
					"00" AFTER 20680 ns,
					"00" AFTER 20700 ns,
					"00" AFTER 20720 ns,
					"00" AFTER 20740 ns,
					"00" AFTER 20760 ns,
					"00" AFTER 20780 ns,
					"00" AFTER 20800 ns,
					"00" AFTER 20820 ns,
					"00" AFTER 20840 ns,
					"00" AFTER 20860 ns,
					"00" AFTER 20880 ns,
					"00" AFTER 20900 ns,
					"00" AFTER 20920 ns,
					"00" AFTER 20940 ns,
					"00" AFTER 20960 ns,
					"00" AFTER 20980 ns,
					"00" AFTER 21000 ns,
					"00" AFTER 21020 ns,
					"00" AFTER 21040 ns,
					"00" AFTER 21060 ns,
					"00" AFTER 21080 ns,
					"00" AFTER 21100 ns,
					"00" AFTER 21120 ns,
					"00" AFTER 21140 ns,
					"00" AFTER 21160 ns,
					"00" AFTER 21180 ns,
					"00" AFTER 21200 ns,
					"00" AFTER 21220 ns,
					"00" AFTER 21240 ns,
					"00" AFTER 21260 ns,
					"00" AFTER 21280 ns,
					"00" AFTER 21300 ns,
					"00" AFTER 21320 ns,
					"00" AFTER 21340 ns,
					"00" AFTER 21360 ns,
					"00" AFTER 21380 ns,
					"00" AFTER 21400 ns,
					"00" AFTER 21420 ns,
					"00" AFTER 21440 ns,
					"00" AFTER 21460 ns,
					"00" AFTER 21480 ns,
					"00" AFTER 21500 ns,
					"00" AFTER 21520 ns,
					"00" AFTER 21540 ns,
					"00" AFTER 21560 ns,
					"00" AFTER 21580 ns,
					"00" AFTER 21600 ns,
					"00" AFTER 21620 ns,
					"00" AFTER 21640 ns,
					"00" AFTER 21660 ns,
					"00" AFTER 21680 ns,
					"00" AFTER 21700 ns,
					"00" AFTER 21720 ns,
					"00" AFTER 21740 ns,
					"00" AFTER 21760 ns,
					"00" AFTER 21780 ns,
					"00" AFTER 21800 ns,
					"00" AFTER 21820 ns,
					"00" AFTER 21840 ns,
					"00" AFTER 21860 ns,
					"00" AFTER 21880 ns,
					"00" AFTER 21900 ns,
					"00" AFTER 21920 ns,
					"00" AFTER 21940 ns,
					"00" AFTER 21960 ns,
					"00" AFTER 21980 ns,
					"00" AFTER 22000 ns,
					"00" AFTER 22020 ns,
					"00" AFTER 22040 ns,
					"00" AFTER 22060 ns,
					"00" AFTER 22080 ns,
					"00" AFTER 22100 ns,
					"00" AFTER 22120 ns,
					"00" AFTER 22140 ns,
					"00" AFTER 22160 ns,
					"00" AFTER 22180 ns,
					"00" AFTER 22200 ns,
					"00" AFTER 22220 ns,
					"00" AFTER 22240 ns,
					"00" AFTER 22260 ns,
					"00" AFTER 22280 ns,
					"00" AFTER 22300 ns,
					"00" AFTER 22320 ns,
					"00" AFTER 22340 ns,
					"00" AFTER 22360 ns,
					"00" AFTER 22380 ns,
					"00" AFTER 22400 ns,
					"00" AFTER 22420 ns,
					"00" AFTER 22440 ns,
					"00" AFTER 22460 ns,
					"00" AFTER 22480 ns,
					"00" AFTER 22500 ns,
					"00" AFTER 22520 ns,
					"00" AFTER 22540 ns,
					"00" AFTER 22560 ns,
					"00" AFTER 22580 ns,
					"00" AFTER 22600 ns,
					"00" AFTER 22620 ns,
					"00" AFTER 22640 ns,
					"00" AFTER 22660 ns,
					"00" AFTER 22680 ns,
					"00" AFTER 22700 ns,
					"00" AFTER 22720 ns,
					"00" AFTER 22740 ns,
					"00" AFTER 22760 ns,
					"00" AFTER 22780 ns,
					"00" AFTER 22800 ns,
					"00" AFTER 22820 ns,
					"00" AFTER 22840 ns,
					"00" AFTER 22860 ns,
					"00" AFTER 22880 ns,
					"00" AFTER 22900 ns,
					"00" AFTER 22920 ns,
					"00" AFTER 22940 ns,
					"00" AFTER 22960 ns,
					"00" AFTER 22980 ns,
					"00" AFTER 23000 ns,
					"00" AFTER 23020 ns,
					"00" AFTER 23040 ns,
					"00" AFTER 23060 ns,
					"00" AFTER 23080 ns,
					"00" AFTER 23100 ns,
					"00" AFTER 23120 ns,
					"00" AFTER 23140 ns,
					"00" AFTER 23160 ns,
					"00" AFTER 23180 ns,
					"00" AFTER 23200 ns,
					"00" AFTER 23220 ns,
					"00" AFTER 23240 ns,
					"00" AFTER 23260 ns,
					"00" AFTER 23280 ns,
					"00" AFTER 23300 ns,
					"00" AFTER 23320 ns,
					"00" AFTER 23340 ns,
					"00" AFTER 23360 ns,
					"00" AFTER 23380 ns,
					"00" AFTER 23400 ns,
					"00" AFTER 23420 ns,
					"00" AFTER 23440 ns,
					"00" AFTER 23460 ns,
					"00" AFTER 23480 ns,
					"00" AFTER 23500 ns,
					"00" AFTER 23520 ns,
					"00" AFTER 23540 ns,
					"00" AFTER 23560 ns,
					"00" AFTER 23580 ns,
					"00" AFTER 23600 ns,
					"00" AFTER 23620 ns,
					"00" AFTER 23640 ns,
					"00" AFTER 23660 ns,
					"00" AFTER 23680 ns,
					"00" AFTER 23700 ns,
					"00" AFTER 23720 ns,
					"00" AFTER 23740 ns,
					"00" AFTER 23760 ns,
					"00" AFTER 23780 ns,
					"00" AFTER 23800 ns,
					"00" AFTER 23820 ns,
					"00" AFTER 23840 ns,
					"00" AFTER 23860 ns,
					"00" AFTER 23880 ns,
					"00" AFTER 23900 ns,
					"00" AFTER 23920 ns,
					"00" AFTER 23940 ns,
					"00" AFTER 23960 ns,
					"00" AFTER 23980 ns,
					"00" AFTER 24000 ns,
					"00" AFTER 24020 ns,
					"00" AFTER 24040 ns,
					"00" AFTER 24060 ns,
					"00" AFTER 24080 ns,
					"00" AFTER 24100 ns,
					"00" AFTER 24120 ns,
					"00" AFTER 24140 ns,
					"00" AFTER 24160 ns,
					"00" AFTER 24180 ns,
					"00" AFTER 24200 ns,
					"00" AFTER 24220 ns,
					"00" AFTER 24240 ns,
					"00" AFTER 24260 ns,
					"00" AFTER 24280 ns,
					"00" AFTER 24300 ns,
					"00" AFTER 24320 ns,
					"00" AFTER 24340 ns,
					"00" AFTER 24360 ns,
					"00" AFTER 24380 ns,
					"00" AFTER 24400 ns,
					"00" AFTER 24420 ns,
					"00" AFTER 24440 ns,
					"00" AFTER 24460 ns,
					"00" AFTER 24480 ns,
					"00" AFTER 24500 ns,
					"00" AFTER 24520 ns,
					"00" AFTER 24540 ns,
					"00" AFTER 24560 ns,
					"00" AFTER 24580 ns,
					"00" AFTER 24600 ns,
					"00" AFTER 24620 ns,
					"00" AFTER 24640 ns,
					"00" AFTER 24660 ns,
					"00" AFTER 24680 ns,
					"00" AFTER 24700 ns,
					"00" AFTER 24720 ns,
					"00" AFTER 24740 ns,
					"00" AFTER 24760 ns,
					"00" AFTER 24780 ns,
					"00" AFTER 24800 ns,
					"00" AFTER 24820 ns,
					"00" AFTER 24840 ns,
					"00" AFTER 24860 ns,
					"00" AFTER 24880 ns,
					"00" AFTER 24900 ns,
					"00" AFTER 24920 ns,
					"00" AFTER 24940 ns,
					"00" AFTER 24960 ns,
					"00" AFTER 24980 ns,
					"00" AFTER 25000 ns,
					"00" AFTER 25020 ns,
					"00" AFTER 25040 ns,
					"00" AFTER 25060 ns,
					"00" AFTER 25080 ns,
					"00" AFTER 25100 ns,
					"00" AFTER 25120 ns,
					"00" AFTER 25140 ns,
					"00" AFTER 25160 ns,
					"00" AFTER 25180 ns,
					"00" AFTER 25200 ns,
					"00" AFTER 25220 ns,
					"00" AFTER 25240 ns,
					"00" AFTER 25260 ns,
					"00" AFTER 25280 ns,
					"00" AFTER 25300 ns,
					"00" AFTER 25320 ns,
					"00" AFTER 25340 ns,
					"00" AFTER 25360 ns,
					"00" AFTER 25380 ns,
					"00" AFTER 25400 ns,
					"00" AFTER 25420 ns,
					"00" AFTER 25440 ns,
					"00" AFTER 25460 ns,
					"00" AFTER 25480 ns,
					"00" AFTER 25500 ns,
					"00" AFTER 25520 ns,
					"00" AFTER 25540 ns,
					"00" AFTER 25560 ns,
					"00" AFTER 25580 ns,
					"00" AFTER 25600 ns,
					"00" AFTER 25620 ns,
					"00" AFTER 25640 ns,
					"00" AFTER 25660 ns,
					"00" AFTER 25680 ns,
					"00" AFTER 25700 ns,
					"00" AFTER 25720 ns,
					"00" AFTER 25740 ns,
					"00" AFTER 25760 ns,
					"00" AFTER 25780 ns,
					"00" AFTER 25800 ns,
					"00" AFTER 25820 ns,
					"00" AFTER 25840 ns,
					"00" AFTER 25860 ns,
					"00" AFTER 25880 ns,
					"00" AFTER 25900 ns,
					"00" AFTER 25920 ns,
					"00" AFTER 25940 ns,
					"00" AFTER 25960 ns,
					"00" AFTER 25980 ns,
					"00" AFTER 26000 ns,
					"00" AFTER 26020 ns,
					"00" AFTER 26040 ns,
					"00" AFTER 26060 ns,
					"00" AFTER 26080 ns,
					"00" AFTER 26100 ns,
					"00" AFTER 26120 ns,
					"00" AFTER 26140 ns,
					"00" AFTER 26160 ns,
					"00" AFTER 26180 ns,
					"00" AFTER 26200 ns,
					"00" AFTER 26220 ns,
					"00" AFTER 26240 ns,
					"00" AFTER 26260 ns,
					"00" AFTER 26280 ns,
					"00" AFTER 26300 ns,
					"00" AFTER 26320 ns,
					"00" AFTER 26340 ns,
					"00" AFTER 26360 ns,
					"00" AFTER 26380 ns,
					"00" AFTER 26400 ns,
					"00" AFTER 26420 ns,
					"00" AFTER 26440 ns,
					"00" AFTER 26460 ns,
					"00" AFTER 26480 ns,
					"00" AFTER 26500 ns,
					"00" AFTER 26520 ns,
					"00" AFTER 26540 ns,
					"00" AFTER 26560 ns,
					"00" AFTER 26580 ns,
					"00" AFTER 26600 ns,
					"00" AFTER 26620 ns,
					"00" AFTER 26640 ns,
					"00" AFTER 26660 ns,
					"00" AFTER 26680 ns,
					"00" AFTER 26700 ns,
					"00" AFTER 26720 ns,
					"00" AFTER 26740 ns,
					"00" AFTER 26760 ns,
					"00" AFTER 26780 ns,
					"00" AFTER 26800 ns,
					"00" AFTER 26820 ns,
					"00" AFTER 26840 ns,
					"00" AFTER 26860 ns,
					"00" AFTER 26880 ns,
					"00" AFTER 26900 ns,
					"00" AFTER 26920 ns,
					"00" AFTER 26940 ns,
					"00" AFTER 26960 ns,
					"00" AFTER 26980 ns,
					"00" AFTER 27000 ns,
					"00" AFTER 27020 ns,
					"00" AFTER 27040 ns,
					"00" AFTER 27060 ns,
					"00" AFTER 27080 ns,
					"00" AFTER 27100 ns,
					"00" AFTER 27120 ns,
					"00" AFTER 27140 ns,
					"00" AFTER 27160 ns,
					"00" AFTER 27180 ns,
					"00" AFTER 27200 ns,
					"00" AFTER 27220 ns,
					"00" AFTER 27240 ns,
					"00" AFTER 27260 ns,
					"00" AFTER 27280 ns,
					"00" AFTER 27300 ns,
					"00" AFTER 27320 ns,
					"00" AFTER 27340 ns,
					"00" AFTER 27360 ns,
					"00" AFTER 27380 ns,
					"00" AFTER 27400 ns,
					"00" AFTER 27420 ns,
					"00" AFTER 27440 ns,
					"00" AFTER 27460 ns,
					"00" AFTER 27480 ns,
					"00" AFTER 27500 ns,
					"00" AFTER 27520 ns,
					"00" AFTER 27540 ns,
					"00" AFTER 27560 ns,
					"00" AFTER 27580 ns,
					"00" AFTER 27600 ns,
					"00" AFTER 27620 ns,
					"00" AFTER 27640 ns,
					"00" AFTER 27660 ns,
					"00" AFTER 27680 ns,
					"00" AFTER 27700 ns,
					"00" AFTER 27720 ns,
					"00" AFTER 27740 ns,
					"00" AFTER 27760 ns,
					"00" AFTER 27780 ns,
					"00" AFTER 27800 ns,
					"00" AFTER 27820 ns,
					"00" AFTER 27840 ns,
					"00" AFTER 27860 ns,
					"00" AFTER 27880 ns,
					"00" AFTER 27900 ns,
					"00" AFTER 27920 ns,
					"00" AFTER 27940 ns,
					"00" AFTER 27960 ns,
					"00" AFTER 27980 ns,
					"00" AFTER 28000 ns,
					"00" AFTER 28020 ns,
					"00" AFTER 28040 ns,
					"00" AFTER 28060 ns,
					"00" AFTER 28080 ns,
					"00" AFTER 28100 ns,
					"00" AFTER 28120 ns,
					"00" AFTER 28140 ns,
					"00" AFTER 28160 ns,
					"00" AFTER 28180 ns,
					"00" AFTER 28200 ns,
					"00" AFTER 28220 ns,
					"01" AFTER 28240 ns,
					"00" AFTER 28260 ns,
					"10" AFTER 28280 ns,
					"00" AFTER 28300 ns,
					"11" AFTER 28320 ns,
					"00" AFTER 28340 ns,
					"00" AFTER 28360 ns,
					"00" AFTER 28380 ns,
					"00" AFTER 28400 ns,
					"00" AFTER 28420 ns,
					"00" AFTER 28440 ns,
					"00" AFTER 28460 ns,
					"00" AFTER 28480 ns,
					"00" AFTER 28500 ns,
					"00" AFTER 28520 ns,
					"00" AFTER 28540 ns,
					"00" AFTER 28560 ns,
					"00" AFTER 28580 ns,
					"00" AFTER 28600 ns,
					"00" AFTER 28620 ns,
					"00" AFTER 28640 ns,
					"00" AFTER 28660 ns,
					"00" AFTER 28680 ns,
					"00" AFTER 28700 ns,
					"00" AFTER 28720 ns,
					"00" AFTER 28740 ns,
					"00" AFTER 28760 ns,
					"00" AFTER 28780 ns,
					"00" AFTER 28800 ns,
					"00" AFTER 28820 ns,
					"00" AFTER 28840 ns,
					"00" AFTER 28860 ns,
					"00" AFTER 28880 ns,
					"00" AFTER 28900 ns,
					"00" AFTER 28920 ns,
					"00" AFTER 28940 ns,
					"00" AFTER 28960 ns,
					"00" AFTER 28980 ns,
					"00" AFTER 29000 ns,
					"00" AFTER 29020 ns,
					"00" AFTER 29040 ns,
					"00" AFTER 29060 ns,
					"00" AFTER 29080 ns,
					"00" AFTER 29100 ns,
					"00" AFTER 29120 ns,
					"00" AFTER 29140 ns,
					"00" AFTER 29160 ns,
					"00" AFTER 29180 ns,
					"00" AFTER 29200 ns,
					"00" AFTER 29220 ns,
					"00" AFTER 29240 ns,
					"00" AFTER 29260 ns,
					"00" AFTER 29280 ns,
					"00" AFTER 29300 ns,
					"00" AFTER 29320 ns,
					"00" AFTER 29340 ns,
					"00" AFTER 29360 ns,
					"00" AFTER 29380 ns,
					"00" AFTER 29400 ns,
					"00" AFTER 29420 ns,
					"00" AFTER 29440 ns,
					"00" AFTER 29460 ns,
					"00" AFTER 29480 ns,
					"00" AFTER 29500 ns,
					"00" AFTER 29520 ns,
					"00" AFTER 29540 ns,
					"00" AFTER 29560 ns,
					"00" AFTER 29580 ns,
					"00" AFTER 29600 ns,
					"00" AFTER 29620 ns,
					"00" AFTER 29640 ns,
					"00" AFTER 29660 ns,
					"00" AFTER 29680 ns,
					"00" AFTER 29700 ns,
					"00" AFTER 29720 ns,
					"00" AFTER 29740 ns,
					"00" AFTER 29760 ns,
					"00" AFTER 29780 ns,
					"00" AFTER 29800 ns,
					"00" AFTER 29820 ns,
					"00" AFTER 29840 ns,
					"00" AFTER 29860 ns,
					"00" AFTER 29880 ns,
					"00" AFTER 29900 ns,
					"00" AFTER 29920 ns,
					"00" AFTER 29940 ns,
					"00" AFTER 29960 ns,
					"00" AFTER 29980 ns,
					"00" AFTER 30000 ns,
					"00" AFTER 30020 ns,
					"00" AFTER 30040 ns,
					"00" AFTER 30060 ns,
					"00" AFTER 30080 ns,
					"00" AFTER 30100 ns,
					"00" AFTER 30120 ns,
					"00" AFTER 30140 ns,
					"00" AFTER 30160 ns,
					"00" AFTER 30180 ns,
					"00" AFTER 30200 ns,
					"00" AFTER 30220 ns,
					"00" AFTER 30240 ns,
					"00" AFTER 30260 ns,
					"00" AFTER 30280 ns,
					"00" AFTER 30300 ns,
					"00" AFTER 30320 ns,
					"00" AFTER 30340 ns,
					"00" AFTER 30360 ns,
					"00" AFTER 30380 ns,
					"00" AFTER 30400 ns,
					"00" AFTER 30420 ns,
					"00" AFTER 30440 ns,
					"00" AFTER 30460 ns,
					"00" AFTER 30480 ns,
					"00" AFTER 30500 ns,
					"00" AFTER 30520 ns,
					"00" AFTER 30540 ns,
					"00" AFTER 30560 ns,
					"00" AFTER 30580 ns,
					"00" AFTER 30600 ns,
					"00" AFTER 30620 ns,
					"00" AFTER 30640 ns,
					"00" AFTER 30660 ns,
					"00" AFTER 30680 ns,
					"00" AFTER 30700 ns,
					"00" AFTER 30720 ns,
					"00" AFTER 30740 ns,
					"00" AFTER 30760 ns,
					"00" AFTER 30780 ns,
					"00" AFTER 30800 ns,
					"00" AFTER 30820 ns,
					"00" AFTER 30840 ns,
					"00" AFTER 30860 ns,
					"00" AFTER 30880 ns,
					"00" AFTER 30900 ns,
					"00" AFTER 30920 ns,
					"00" AFTER 30940 ns,
					"00" AFTER 30960 ns;

ControlRegisters <=  "000000000000000000000000000" AFTER 00020 ns,
							"000000000000000000000000001" AFTER 00040 ns,
							"000000000000000000000000000" AFTER 00060 ns,
							"000000000000000000000000001" AFTER 00080 ns,
							"000000000000000000000000000" AFTER 00100 ns,
							"000000000000000000000000001" AFTER 00120 ns,
							"000000000000000000000000000" AFTER 00140 ns,
							"000000000000000000000000001" AFTER 00160 ns,
							"000000000000000000000000000" AFTER 00180 ns,
							"000000000000000000000000001" AFTER 00200 ns,
							"000000000000000000000000000" AFTER 00220 ns,
							"000000000000000000000000001" AFTER 00240 ns,
							"000000000000000000000000000" AFTER 00260 ns,
							"000000000000000000000000001" AFTER 00280 ns,
							"000000000000000000000000000" AFTER 00300 ns,
							"000000000000000000000000001" AFTER 00320 ns,
							"000000000000000000000000000" AFTER 00340 ns,
							"000000000000000000000000001" AFTER 00360 ns,
							"000000000000000000000000000" AFTER 00380 ns,
							"000000000000000000000000001" AFTER 00400 ns,
							"000000000000000000000000000" AFTER 00420 ns,
							"000000000000000000000000001" AFTER 00440 ns,
							"000000000000000000000000000" AFTER 00460 ns,
							"000000000000000000000000001" AFTER 00480 ns,
							"000000000000000000000000000" AFTER 00500 ns,
							"000000000000000000000000001" AFTER 00520 ns,
							"000000000000000000000000000" AFTER 00540 ns,
							"000000000000000000000000001" AFTER 00560 ns,
							"000000000000000000000000000" AFTER 00580 ns,
							"000000000000000000000000001" AFTER 00600 ns,
							"000000000000000000000000000" AFTER 00620 ns,
							"000000000000000000000000001" AFTER 00640 ns,
							"000000000000000000000000000" AFTER 00660 ns,
							"000000000000000000000000001" AFTER 00680 ns,
							"000000000000000000000000000" AFTER 00700 ns,
							"000000000000000000000000001" AFTER 00720 ns,
							"000000000000000000000000000" AFTER 00740 ns,
							"000000000000000000000000001" AFTER 00760 ns,
							"000000000000000000000000000" AFTER 00780 ns,
							"000000000000000000000000001" AFTER 00800 ns,
							"000000000000000000000000000" AFTER 00820 ns,
							"000000000000000000000000001" AFTER 00840 ns,
							"000000000000000000000000000" AFTER 00860 ns,
							"000000000000000000000000001" AFTER 00880 ns,
							"000000000000000000000000000" AFTER 00900 ns,
							"000000000000000000000000001" AFTER 00920 ns,
							"000000000000000000000000000" AFTER 00940 ns,
							"000000000000000000000000001" AFTER 00960 ns,
							"000000000000000000000000000" AFTER 00980 ns,
							"000000000000000000000000001" AFTER 01000 ns,
							"000000000000000000000000000" AFTER 01020 ns,
							"000000000000000000000000001" AFTER 01040 ns,
							"000000000000000000000000000" AFTER 01060 ns,
							"000000000000000000000000001" AFTER 01080 ns,
							"000000000000000000000000000" AFTER 01100 ns,
							"000000000000000000000000001" AFTER 01120 ns,
							"000000000000000000000000000" AFTER 01140 ns,
							"000000000000000000000000001" AFTER 01160 ns,
							"000000000000000000000000000" AFTER 01180 ns,
							"000000000000000000000000001" AFTER 01200 ns,
							"000000000000000000000000000" AFTER 01220 ns,
							"000000000000000000000000001" AFTER 01240 ns,
							"000000000000000000000000000" AFTER 01260 ns,
							"000000000000000000000000001" AFTER 01280 ns,
							"000000000000000000000000000" AFTER 01300 ns,
							"000000000000000000000000010" AFTER 01320 ns,
							"000000000000000000000000000" AFTER 01340 ns,
							"000000000000000000000000010" AFTER 01360 ns,
							"000000000000000000000000000" AFTER 01380 ns,
							"000000000000000000000000010" AFTER 01400 ns,
							"000000000000000000000000000" AFTER 01420 ns,
							"000000000000000000000000010" AFTER 01440 ns,
							"000000000000000000000000000" AFTER 01460 ns,
							"000000000000000000000000010" AFTER 01480 ns,
							"000000000000000000000000000" AFTER 01500 ns,
							"000000000000000000000000010" AFTER 01520 ns,
							"000000000000000000000000000" AFTER 01540 ns,
							"000000000000000000000000010" AFTER 01560 ns,
							"000000000000000000000000000" AFTER 01580 ns,
							"000000000000000000000000010" AFTER 01600 ns,
							"000000000000000000000000000" AFTER 01620 ns,
							"000000000000000000000000010" AFTER 01640 ns,
							"000000000000000000000000000" AFTER 01660 ns,
							"000000000000000000000000010" AFTER 01680 ns,
							"000000000000000000000000000" AFTER 01700 ns,
							"000000000000000000000000010" AFTER 01720 ns,
							"000000000000000000000000000" AFTER 01740 ns,
							"000000000000000000000000010" AFTER 01760 ns,
							"000000000000000000000000000" AFTER 01780 ns,
							"000000000000000000000000010" AFTER 01800 ns,
							"000000000000000000000000000" AFTER 01820 ns,
							"000000000000000000000000010" AFTER 01840 ns,
							"000000000000000000000000000" AFTER 01860 ns,
							"000000000000000000000000010" AFTER 01880 ns,
							"000000000000000000000000000" AFTER 01900 ns,
							"000000000000000000000000010" AFTER 01920 ns,
							"000000000000000000000000000" AFTER 01940 ns,
							"000000000000000000000000010" AFTER 01960 ns,
							"000000000000000000000000000" AFTER 01980 ns,
							"000000000000000000000000010" AFTER 02000 ns,
							"000000000000000000000000000" AFTER 02020 ns,
							"000000000000000000000000010" AFTER 02040 ns,
							"000000000000000000000000000" AFTER 02060 ns,
							"000000000000000000000000010" AFTER 02080 ns,
							"000000000000000000000000000" AFTER 02100 ns,
							"000000000000000000000000010" AFTER 02120 ns,
							"000000000000000000000000000" AFTER 02140 ns,
							"000000000000000000000000010" AFTER 02160 ns,
							"000000000000000000000000000" AFTER 02180 ns,
							"000000000000000000000000010" AFTER 02200 ns,
							"000000000000000000000000000" AFTER 02220 ns,
							"000000000000000000000000010" AFTER 02240 ns,
							"000000000000000000000000000" AFTER 02260 ns,
							"000000000000000000000000010" AFTER 02280 ns,
							"000000000000000000000000000" AFTER 02300 ns,
							"000000000000000000000000010" AFTER 02320 ns,
							"000000000000000000000000000" AFTER 02340 ns,
							"000000000000000000000000010" AFTER 02360 ns,
							"000000000000000000000000000" AFTER 02380 ns,
							"000000000000000000000000010" AFTER 02400 ns,
							"000000000000000000000000000" AFTER 02420 ns,
							"000000000000000000000000010" AFTER 02440 ns,
							"000000000000000000000000000" AFTER 02460 ns,
							"000000000000000000000000010" AFTER 02480 ns,
							"000000000000000000000000000" AFTER 02500 ns,
							"000000000000000000000000010" AFTER 02520 ns,
							"000000000000000000000000000" AFTER 02540 ns,
							"000000000000000000000000010" AFTER 02560 ns,
							"000000000000000000000000000" AFTER 02580 ns,
							"000000000000000000000000100" AFTER 02600 ns,
							"000000000000000000000000000" AFTER 02620 ns,
							"000000000000000000000000100" AFTER 02640 ns,
							"000000000000000000000000000" AFTER 02660 ns,
							"000000000000000000000000100" AFTER 02680 ns,
							"000000000000000000000000000" AFTER 02700 ns,
							"000000000000000000000000100" AFTER 02720 ns,
							"000000000000000000000000000" AFTER 02740 ns,
							"000000000000000000000000100" AFTER 02760 ns,
							"000000000000000000000000000" AFTER 02780 ns,
							"000000000000000000000000100" AFTER 02800 ns,
							"000000000000000000000000000" AFTER 02820 ns,
							"000000000000000000000000100" AFTER 02840 ns,
							"000000000000000000000000000" AFTER 02860 ns,
							"000000000000000000000000100" AFTER 02880 ns,
							"000000000000000000000000000" AFTER 02900 ns,
							"000000000000000000000000100" AFTER 02920 ns,
							"000000000000000000000000000" AFTER 02940 ns,
							"000000000000000000000000100" AFTER 02960 ns,
							"000000000000000000000000000" AFTER 02980 ns,
							"000000000000000000000000100" AFTER 03000 ns,
							"000000000000000000000000000" AFTER 03020 ns,
							"000000000000000000000000100" AFTER 03040 ns,
							"000000000000000000000000000" AFTER 03060 ns,
							"000000000000000000000000100" AFTER 03080 ns,
							"000000000000000000000000000" AFTER 03100 ns,
							"000000000000000000000000100" AFTER 03120 ns,
							"000000000000000000000000000" AFTER 03140 ns,
							"000000000000000000000000100" AFTER 03160 ns,
							"000000000000000000000000000" AFTER 03180 ns,
							"000000000000000000000000100" AFTER 03200 ns,
							"000000000000000000000000000" AFTER 03220 ns,
							"000000000000000000000000100" AFTER 03240 ns,
							"000000000000000000000000000" AFTER 03260 ns,
							"000000000000000000000000100" AFTER 03280 ns,
							"000000000000000000000000000" AFTER 03300 ns,
							"000000000000000000000000100" AFTER 03320 ns,
							"000000000000000000000000000" AFTER 03340 ns,
							"000000000000000000000000100" AFTER 03360 ns,
							"000000000000000000000000000" AFTER 03380 ns,
							"000000000000000000000000100" AFTER 03400 ns,
							"000000000000000000000000000" AFTER 03420 ns,
							"000000000000000000000000100" AFTER 03440 ns,
							"000000000000000000000000000" AFTER 03460 ns,
							"000000000000000000000000100" AFTER 03480 ns,
							"000000000000000000000000000" AFTER 03500 ns,
							"000000000000000000000000100" AFTER 03520 ns,
							"000000000000000000000000000" AFTER 03540 ns,
							"000000000000000000000000100" AFTER 03560 ns,
							"000000000000000000000000000" AFTER 03580 ns,
							"000000000000000000000000100" AFTER 03600 ns,
							"000000000000000000000000000" AFTER 03620 ns,
							"000000000000000000000000100" AFTER 03640 ns,
							"000000000000000000000000000" AFTER 03660 ns,
							"000000000000000000000000100" AFTER 03680 ns,
							"000000000000000000000000000" AFTER 03700 ns,
							"000000000000000000000000100" AFTER 03720 ns,
							"000000000000000000000000000" AFTER 03740 ns,
							"000000000000000000000000100" AFTER 03760 ns,
							"000000000000000000000000000" AFTER 03780 ns,
							"000000000000000000000000100" AFTER 03800 ns,
							"000000000000000000000000000" AFTER 03820 ns,
							"000000000000000000000000100" AFTER 03840 ns,
							"000000000000000000000000000" AFTER 03860 ns,
							"000000000000000000000001000" AFTER 03880 ns,
							"000000000000000000000000000" AFTER 03900 ns,
							"000000000000000000000001000" AFTER 03920 ns,
							"000000000000000000000000000" AFTER 03940 ns,
							"000000000000000000000001000" AFTER 03960 ns,
							"000000000000000000000000000" AFTER 03980 ns,
							"000000000000000000000001000" AFTER 04000 ns,
							"000000000000000000000000000" AFTER 04020 ns,
							"000000000000000000000001000" AFTER 04040 ns,
							"000000000000000000000000000" AFTER 04060 ns,
							"000000000000000000000001000" AFTER 04080 ns,
							"000000000000000000000000000" AFTER 04100 ns,
							"000000000000000000000001000" AFTER 04120 ns,
							"000000000000000000000000000" AFTER 04140 ns,
							"000000000000000000000001000" AFTER 04160 ns,
							"000000000000000000000000000" AFTER 04180 ns,
							"000000000000000000000001000" AFTER 04200 ns,
							"000000000000000000000000000" AFTER 04220 ns,
							"000000000000000000000001000" AFTER 04240 ns,
							"000000000000000000000000000" AFTER 04260 ns,
							"000000000000000000000001000" AFTER 04280 ns,
							"000000000000000000000000000" AFTER 04300 ns,
							"000000000000000000000001000" AFTER 04320 ns,
							"000000000000000000000000000" AFTER 04340 ns,
							"000000000000000000000001000" AFTER 04360 ns,
							"000000000000000000000000000" AFTER 04380 ns,
							"000000000000000000000001000" AFTER 04400 ns,
							"000000000000000000000000000" AFTER 04420 ns,
							"000000000000000000000001000" AFTER 04440 ns,
							"000000000000000000000000000" AFTER 04460 ns,
							"000000000000000000000001000" AFTER 04480 ns,
							"000000000000000000000000000" AFTER 04500 ns,
							"000000000000000000000001000" AFTER 04520 ns,
							"000000000000000000000000000" AFTER 04540 ns,
							"000000000000000000000001000" AFTER 04560 ns,
							"000000000000000000000000000" AFTER 04580 ns,
							"000000000000000000000001000" AFTER 04600 ns,
							"000000000000000000000000000" AFTER 04620 ns,
							"000000000000000000000001000" AFTER 04640 ns,
							"000000000000000000000000000" AFTER 04660 ns,
							"000000000000000000000001000" AFTER 04680 ns,
							"000000000000000000000000000" AFTER 04700 ns,
							"000000000000000000000001000" AFTER 04720 ns,
							"000000000000000000000000000" AFTER 04740 ns,
							"000000000000000000000001000" AFTER 04760 ns,
							"000000000000000000000000000" AFTER 04780 ns,
							"000000000000000000000001000" AFTER 04800 ns,
							"000000000000000000000000000" AFTER 04820 ns,
							"000000000000000000000001000" AFTER 04840 ns,
							"000000000000000000000000000" AFTER 04860 ns,
							"000000000000000000000001000" AFTER 04880 ns,
							"000000000000000000000000000" AFTER 04900 ns,
							"000000000000000000000001000" AFTER 04920 ns,
							"000000000000000000000000000" AFTER 04940 ns,
							"000000000000000000000001000" AFTER 04960 ns,
							"000000000000000000000000000" AFTER 04980 ns,
							"000000000000000000000001000" AFTER 05000 ns,
							"000000000000000000000000000" AFTER 05020 ns,
							"000000000000000000000001000" AFTER 05040 ns,
							"000000000000000000000000000" AFTER 05060 ns,
							"000000000000000000000001000" AFTER 05080 ns,
							"000000000000000000000000000" AFTER 05100 ns,
							"000000000000000000000001000" AFTER 05120 ns,
							"000000000000000000000000000" AFTER 05140 ns,
							"000000000000000000000100000" AFTER 05160 ns,
							"000000000000000000000000000" AFTER 05180 ns,
							"000000000000000000000100000" AFTER 05200 ns,
							"000000000000000000000000000" AFTER 05220 ns,
							"000000000000000000000100000" AFTER 05240 ns,
							"000000000000000000000000000" AFTER 05260 ns,
							"000000000000000000000100000" AFTER 05280 ns,
							"000000000000000000000000000" AFTER 05300 ns,
							"000000000000000000000100000" AFTER 05320 ns,
							"000000000000000000000000000" AFTER 05340 ns,
							"000000000000000000000100000" AFTER 05360 ns,
							"000000000000000000000000000" AFTER 05380 ns,
							"000000000000000000000100000" AFTER 05400 ns,
							"000000000000000000000000000" AFTER 05420 ns,
							"000000000000000000000100000" AFTER 05440 ns,
							"000000000000000000000000000" AFTER 05460 ns,
							"000000000000000000000100000" AFTER 05480 ns,
							"000000000000000000000000000" AFTER 05500 ns,
							"000000000000000000000100000" AFTER 05520 ns,
							"000000000000000000000000000" AFTER 05540 ns,
							"000000000000000000000100000" AFTER 05560 ns,
							"000000000000000000000000000" AFTER 05580 ns,
							"000000000000000000000100000" AFTER 05600 ns,
							"000000000000000000000000000" AFTER 05620 ns,
							"000000000000000000000100000" AFTER 05640 ns,
							"000000000000000000000000000" AFTER 05660 ns,
							"000000000000000000000100000" AFTER 05680 ns,
							"000000000000000000000000000" AFTER 05700 ns,
							"000000000000000000000100000" AFTER 05720 ns,
							"000000000000000000000000000" AFTER 05740 ns,
							"000000000000000000000100000" AFTER 05760 ns,
							"000000000000000000000000000" AFTER 05780 ns,
							"000000000000000000000100000" AFTER 05800 ns,
							"000000000000000000000000000" AFTER 05820 ns,
							"000000000000000000000100000" AFTER 05840 ns,
							"000000000000000000000000000" AFTER 05860 ns,
							"000000000000000000000100000" AFTER 05880 ns,
							"000000000000000000000000000" AFTER 05900 ns,
							"000000000000000000000100000" AFTER 05920 ns,
							"000000000000000000000000000" AFTER 05940 ns,
							"000000000000000000000100000" AFTER 05960 ns,
							"000000000000000000000000000" AFTER 05980 ns,
							"000000000000000000000100000" AFTER 06000 ns,
							"000000000000000000000000000" AFTER 06020 ns,
							"000000000000000000000100000" AFTER 06040 ns,
							"000000000000000000000000000" AFTER 06060 ns,
							"000000000000000000000100000" AFTER 06080 ns,
							"000000000000000000000000000" AFTER 06100 ns,
							"000000000000000000000100000" AFTER 06120 ns,
							"000000000000000000000000000" AFTER 06140 ns,
							"000000000000000000000100000" AFTER 06160 ns,
							"000000000000000000000000000" AFTER 06180 ns,
							"000000000000000000000100000" AFTER 06200 ns,
							"000000000000000000000000000" AFTER 06220 ns,
							"000000000000000000000100000" AFTER 06240 ns,
							"000000000000000000000000000" AFTER 06260 ns,
							"000000000000000000000100000" AFTER 06280 ns,
							"000000000000000000000000000" AFTER 06300 ns,
							"000000000000000000000100000" AFTER 06320 ns,
							"000000000000000000000000000" AFTER 06340 ns,
							"000000000000000000000100000" AFTER 06360 ns,
							"000000000000000000000000000" AFTER 06380 ns,
							"000000000000000000000100000" AFTER 06400 ns,
							"000000000000000000000000000" AFTER 06420 ns,
							"000000000000000000000010000" AFTER 06440 ns,
							"000000000000000000000000000" AFTER 06460 ns,
							"000000000000000000000010000" AFTER 06480 ns,
							"000000000000000000000000000" AFTER 06500 ns,
							"000000000000000000000010000" AFTER 06520 ns,
							"000000000000000000000000000" AFTER 06540 ns,
							"000000000000000000000010000" AFTER 06560 ns,
							"000000000000000000000000000" AFTER 06580 ns,
							"000000000000000000000010000" AFTER 06600 ns,
							"000000000000000000000000000" AFTER 06620 ns,
							"000000000000000000000010000" AFTER 06640 ns,
							"000000000000000000000000000" AFTER 06660 ns,
							"000000000000000000000010000" AFTER 06680 ns,
							"000000000000000000000000000" AFTER 06700 ns,
							"000000000000000000000010000" AFTER 06720 ns,
							"000000000000000000000000000" AFTER 06740 ns,
							"000000000000000000000010000" AFTER 06760 ns,
							"000000000000000000000000000" AFTER 06780 ns,
							"000000000000000000000010000" AFTER 06800 ns,
							"000000000000000000000000000" AFTER 06820 ns,
							"000000000000000000000010000" AFTER 06840 ns,
							"000000000000000000000000000" AFTER 06860 ns,
							"000000000000000000000010000" AFTER 06880 ns,
							"000000000000000000000000000" AFTER 06900 ns,
							"000000000000000000000010000" AFTER 06920 ns,
							"000000000000000000000000000" AFTER 06940 ns,
							"000000000000000000000010000" AFTER 06960 ns,
							"000000000000000000000000000" AFTER 06980 ns,
							"000000000000000000000010000" AFTER 07000 ns,
							"000000000000000000000000000" AFTER 07020 ns,
							"000000000000000000000010000" AFTER 07040 ns,
							"000000000000000000000000000" AFTER 07060 ns,
							"000000000000000000000010000" AFTER 07080 ns,
							"000000000000000000000000000" AFTER 07100 ns,
							"000000000000000000000010000" AFTER 07120 ns,
							"000000000000000000000000000" AFTER 07140 ns,
							"000000000000000000000010000" AFTER 07160 ns,
							"000000000000000000000000000" AFTER 07180 ns,
							"000000000000000000000010000" AFTER 07200 ns,
							"000000000000000000000000000" AFTER 07220 ns,
							"000000000000000000000010000" AFTER 07240 ns,
							"000000000000000000000000000" AFTER 07260 ns,
							"000000000000000000000010000" AFTER 07280 ns,
							"000000000000000000000000000" AFTER 07300 ns,
							"000000000000000000000010000" AFTER 07320 ns,
							"000000000000000000000000000" AFTER 07340 ns,
							"000000000000000000000010000" AFTER 07360 ns,
							"000000000000000000000000000" AFTER 07380 ns,
							"000000000000000000000010000" AFTER 07400 ns,
							"000000000000000000000000000" AFTER 07420 ns,
							"000000000000000000000010000" AFTER 07440 ns,
							"000000000000000000000000000" AFTER 07460 ns,
							"000000000000000000000010000" AFTER 07480 ns,
							"000000000000000000000000000" AFTER 07500 ns,
							"000000000000000000000010000" AFTER 07520 ns,
							"000000000000000000000000000" AFTER 07540 ns,
							"000000000000000000000010000" AFTER 07560 ns,
							"000000000000000000000000000" AFTER 07580 ns,
							"000000000000000000000010000" AFTER 07600 ns,
							"000000000000000000000000000" AFTER 07620 ns,
							"000000000000000000000010000" AFTER 07640 ns,
							"000000000000000000000000000" AFTER 07660 ns,
							"000000000000000000000010000" AFTER 07680 ns,
							"000000000000000000000000000" AFTER 07700 ns,
							"000000000000000000001000000" AFTER 07720 ns,
							"000000000000000000000000000" AFTER 07740 ns,
							"000000000000000000001000000" AFTER 07760 ns,
							"000000000000000000000000000" AFTER 07780 ns,
							"000000000000000000001000000" AFTER 07800 ns,
							"000000000000000000000000000" AFTER 07820 ns,
							"000000000000000000001000000" AFTER 07840 ns,
							"000000000000000000000000000" AFTER 07860 ns,
							"000000000000000000001000000" AFTER 07880 ns,
							"000000000000000000000000000" AFTER 07900 ns,
							"000000000000000000001000000" AFTER 07920 ns,
							"000000000000000000000000000" AFTER 07940 ns,
							"000000000000000000001000000" AFTER 07960 ns,
							"000000000000000000000000000" AFTER 07980 ns,
							"000000000000000000001000000" AFTER 08000 ns,
							"000000000000000000000000000" AFTER 08020 ns,
							"000000000000000000001000000" AFTER 08040 ns,
							"000000000000000000000000000" AFTER 08060 ns,
							"000000000000000000001000000" AFTER 08080 ns,
							"000000000000000000000000000" AFTER 08100 ns,
							"000000000000000000001000000" AFTER 08120 ns,
							"000000000000000000000000000" AFTER 08140 ns,
							"000000000000000000001000000" AFTER 08160 ns,
							"000000000000000000000000000" AFTER 08180 ns,
							"000000000000000000001000000" AFTER 08200 ns,
							"000000000000000000000000000" AFTER 08220 ns,
							"000000000000000000001000000" AFTER 08240 ns,
							"000000000000000000000000000" AFTER 08260 ns,
							"000000000000000000001000000" AFTER 08280 ns,
							"000000000000000000000000000" AFTER 08300 ns,
							"000000000000000000001000000" AFTER 08320 ns,
							"000000000000000000000000000" AFTER 08340 ns,
							"000000000000000000001000000" AFTER 08360 ns,
							"000000000000000000000000000" AFTER 08380 ns,
							"000000000000000000001000000" AFTER 08400 ns,
							"000000000000000000000000000" AFTER 08420 ns,
							"000000000000000000001000000" AFTER 08440 ns,
							"000000000000000000000000000" AFTER 08460 ns,
							"000000000000000000001000000" AFTER 08480 ns,
							"000000000000000000000000000" AFTER 08500 ns,
							"000000000000000000001000000" AFTER 08520 ns,
							"000000000000000000000000000" AFTER 08540 ns,
							"000000000000000000001000000" AFTER 08560 ns,
							"000000000000000000000000000" AFTER 08580 ns,
							"000000000000000000001000000" AFTER 08600 ns,
							"000000000000000000000000000" AFTER 08620 ns,
							"000000000000000000001000000" AFTER 08640 ns,
							"000000000000000000000000000" AFTER 08660 ns,
							"000000000000000000001000000" AFTER 08680 ns,
							"000000000000000000000000000" AFTER 08700 ns,
							"000000000000000000001000000" AFTER 08720 ns,
							"000000000000000000000000000" AFTER 08740 ns,
							"000000000000000000001000000" AFTER 08760 ns,
							"000000000000000000000000000" AFTER 08780 ns,
							"000000000000000000001000000" AFTER 08800 ns,
							"000000000000000000000000000" AFTER 08820 ns,
							"000000000000000000001000000" AFTER 08840 ns,
							"000000000000000000000000000" AFTER 08860 ns,
							"000000000000000000001000000" AFTER 08880 ns,
							"000000000000000000000000000" AFTER 08900 ns,
							"000000000000000000001000000" AFTER 08920 ns,
							"000000000000000000000000000" AFTER 08940 ns,
							"000000000000000000001000000" AFTER 08960 ns,
							"000000000000000000000000000" AFTER 08980 ns,
							"000000000000000000010000000" AFTER 09000 ns,
							"000000000000000000000000000" AFTER 09020 ns,
							"000000000000000000010000000" AFTER 09040 ns,
							"000000000000000000000000000" AFTER 09060 ns,
							"000000000000000000010000000" AFTER 09080 ns,
							"000000000000000000000000000" AFTER 09100 ns,
							"000000000000000000010000000" AFTER 09120 ns,
							"000000000000000000000000000" AFTER 09140 ns,
							"000000000000000000010000000" AFTER 09160 ns,
							"000000000000000000000000000" AFTER 09180 ns,
							"000000000000000000010000000" AFTER 09200 ns,
							"000000000000000000000000000" AFTER 09220 ns,
							"000000000000000000010000000" AFTER 09240 ns,
							"000000000000000000000000000" AFTER 09260 ns,
							"000000000000000000010000000" AFTER 09280 ns,
							"000000000000000000000000000" AFTER 09300 ns,
							"000000000000000000010000000" AFTER 09320 ns,
							"000000000000000000000000000" AFTER 09340 ns,
							"000000000000000000010000000" AFTER 09360 ns,
							"000000000000000000000000000" AFTER 09380 ns,
							"000000000000000000010000000" AFTER 09400 ns,
							"000000000000000000000000000" AFTER 09420 ns,
							"000000000000000000010000000" AFTER 09440 ns,
							"000000000000000000000000000" AFTER 09460 ns,
							"000000000000000000010000000" AFTER 09480 ns,
							"000000000000000000000000000" AFTER 09500 ns,
							"000000000000000000010000000" AFTER 09520 ns,
							"000000000000000000000000000" AFTER 09540 ns,
							"000000000000000000010000000" AFTER 09560 ns,
							"000000000000000000000000000" AFTER 09580 ns,
							"000000000000000000010000000" AFTER 09600 ns,
							"000000000000000000000000000" AFTER 09620 ns,
							"000000000000000000010000000" AFTER 09640 ns,
							"000000000000000000000000000" AFTER 09660 ns,
							"000000000000000000010000000" AFTER 09680 ns,
							"000000000000000000000000000" AFTER 09700 ns,
							"000000000000000000010000000" AFTER 09720 ns,
							"000000000000000000000000000" AFTER 09740 ns,
							"000000000000000000010000000" AFTER 09760 ns,
							"000000000000000000000000000" AFTER 09780 ns,
							"000000000000000000010000000" AFTER 09800 ns,
							"000000000000000000000000000" AFTER 09820 ns,
							"000000000000000000010000000" AFTER 09840 ns,
							"000000000000000000000000000" AFTER 09860 ns,
							"000000000000000000010000000" AFTER 09880 ns,
							"000000000000000000000000000" AFTER 09900 ns,
							"000000000000000000010000000" AFTER 09920 ns,
							"000000000000000000000000000" AFTER 09940 ns,
							"000000000000000000010000000" AFTER 09960 ns,
							"000000000000000000000000000" AFTER 09980 ns,
							"000000000000000000010000000" AFTER 10000 ns,
							"000000000000000000000000000" AFTER 10020 ns,
							"000000000000000000010000000" AFTER 10040 ns,
							"000000000000000000000000000" AFTER 10060 ns,
							"000000000000000000010000000" AFTER 10080 ns,
							"000000000000000000000000000" AFTER 10100 ns,
							"000000000000000000010000000" AFTER 10120 ns,
							"000000000000000000000000000" AFTER 10140 ns,
							"000000000000000000010000000" AFTER 10160 ns,
							"000000000000000000000000000" AFTER 10180 ns,
							"000000000000000000010000000" AFTER 10200 ns,
							"000000000000000000000000000" AFTER 10220 ns,
							"000000000000000000010000000" AFTER 10240 ns,
							"000000000000000000000000000" AFTER 10260 ns,
							"000000000000000000100000000" AFTER 10280 ns,
							"000000000000000000000000000" AFTER 10300 ns,
							"000000000000000000100000000" AFTER 10320 ns,
							"000000000000000000000000000" AFTER 10340 ns,
							"000000000000000000100000000" AFTER 10360 ns,
							"000000000000000000000000000" AFTER 10380 ns,
							"000000000000000000100000000" AFTER 10400 ns,
							"000000000000000000000000000" AFTER 10420 ns,
							"000000000000000000100000000" AFTER 10440 ns,
							"000000000000000000000000000" AFTER 10460 ns,
							"000000000000000000100000000" AFTER 10480 ns,
							"000000000000000000000000000" AFTER 10500 ns,
							"000000000000000000100000000" AFTER 10520 ns,
							"000000000000000000000000000" AFTER 10540 ns,
							"000000000000000000100000000" AFTER 10560 ns,
							"000000000000000000000000000" AFTER 10580 ns,
							"000000000000000000100000000" AFTER 10600 ns,
							"000000000000000000000000000" AFTER 10620 ns,
							"000000000000000000100000000" AFTER 10640 ns,
							"000000000000000000000000000" AFTER 10660 ns,
							"000000000000000000100000000" AFTER 10680 ns,
							"000000000000000000000000000" AFTER 10700 ns,
							"000000000000000000100000000" AFTER 10720 ns,
							"000000000000000000000000000" AFTER 10740 ns,
							"000000000000000000100000000" AFTER 10760 ns,
							"000000000000000000000000000" AFTER 10780 ns,
							"000000000000000000100000000" AFTER 10800 ns,
							"000000000000000000000000000" AFTER 10820 ns,
							"000000000000000000100000000" AFTER 10840 ns,
							"000000000000000000000000000" AFTER 10860 ns,
							"000000000000000000100000000" AFTER 10880 ns,
							"000000000000000000000000000" AFTER 10900 ns,
							"000000000000000000100000000" AFTER 10920 ns,
							"000000000000000000000000000" AFTER 10940 ns,
							"000000000000000000100000000" AFTER 10960 ns,
							"000000000000000000000000000" AFTER 10980 ns,
							"000000000000000000100000000" AFTER 11000 ns,
							"000000000000000000000000000" AFTER 11020 ns,
							"000000000000000000100000000" AFTER 11040 ns,
							"000000000000000000000000000" AFTER 11060 ns,
							"000000000000000000100000000" AFTER 11080 ns,
							"000000000000000000000000000" AFTER 11100 ns,
							"000000000000000000100000000" AFTER 11120 ns,
							"000000000000000000000000000" AFTER 11140 ns,
							"000000000000000000100000000" AFTER 11160 ns,
							"000000000000000000000000000" AFTER 11180 ns,
							"000000000000000000100000000" AFTER 11200 ns,
							"000000000000000000000000000" AFTER 11220 ns,
							"000000000000000000100000000" AFTER 11240 ns,
							"000000000000000000000000000" AFTER 11260 ns,
							"000000000000000000100000000" AFTER 11280 ns,
							"000000000000000000000000000" AFTER 11300 ns,
							"000000000000000000100000000" AFTER 11320 ns,
							"000000000000000000000000000" AFTER 11340 ns,
							"000000000000000000100000000" AFTER 11360 ns,
							"000000000000000000000000000" AFTER 11380 ns,
							"000000000000000000100000000" AFTER 11400 ns,
							"000000000000000000000000000" AFTER 11420 ns,
							"000000000000000000100000000" AFTER 11440 ns,
							"000000000000000000000000000" AFTER 11460 ns,
							"000000000000000000100000000" AFTER 11480 ns,
							"000000000000000000000000000" AFTER 11500 ns,
							"000000000000000000100000000" AFTER 11520 ns,
							"000000000000000000000000000" AFTER 11540 ns,
							"000000000000000001000000000" AFTER 11560 ns,
							"000000000000000000000000000" AFTER 11580 ns,
							"000000000000000001000000000" AFTER 11600 ns,
							"000000000000000000000000000" AFTER 11620 ns,
							"000000000000000001000000000" AFTER 11640 ns,
							"000000000000000000000000000" AFTER 11660 ns,
							"000000000000000001000000000" AFTER 11680 ns,
							"000000000000000000000000000" AFTER 11700 ns,
							"000000000000000001000000000" AFTER 11720 ns,
							"000000000000000000000000000" AFTER 11740 ns,
							"000000000000000001000000000" AFTER 11760 ns,
							"000000000000000000000000000" AFTER 11780 ns,
							"000000000000000001000000000" AFTER 11800 ns,
							"000000000000000000000000000" AFTER 11820 ns,
							"000000000000000001000000000" AFTER 11840 ns,
							"000000000000000000000000000" AFTER 11860 ns,
							"000000000000000001000000000" AFTER 11880 ns,
							"000000000000000000000000000" AFTER 11900 ns,
							"000000000000000001000000000" AFTER 11920 ns,
							"000000000000000000000000000" AFTER 11940 ns,
							"000000000000000001000000000" AFTER 11960 ns,
							"000000000000000000000000000" AFTER 11980 ns,
							"000000000000000001000000000" AFTER 12000 ns,
							"000000000000000000000000000" AFTER 12020 ns,
							"000000000000000001000000000" AFTER 12040 ns,
							"000000000000000000000000000" AFTER 12060 ns,
							"000000000000000001000000000" AFTER 12080 ns,
							"000000000000000000000000000" AFTER 12100 ns,
							"000000000000000001000000000" AFTER 12120 ns,
							"000000000000000000000000000" AFTER 12140 ns,
							"000000000000000001000000000" AFTER 12160 ns,
							"000000000000000000000000000" AFTER 12180 ns,
							"000000000000000001000000000" AFTER 12200 ns,
							"000000000000000000000000000" AFTER 12220 ns,
							"000000000000000001000000000" AFTER 12240 ns,
							"000000000000000000000000000" AFTER 12260 ns,
							"000000000000000001000000000" AFTER 12280 ns,
							"000000000000000000000000000" AFTER 12300 ns,
							"000000000000000001000000000" AFTER 12320 ns,
							"000000000000000000000000000" AFTER 12340 ns,
							"000000000000000001000000000" AFTER 12360 ns,
							"000000000000000000000000000" AFTER 12380 ns,
							"000000000000000001000000000" AFTER 12400 ns,
							"000000000000000000000000000" AFTER 12420 ns,
							"000000000000000001000000000" AFTER 12440 ns,
							"000000000000000000000000000" AFTER 12460 ns,
							"000000000000000001000000000" AFTER 12480 ns,
							"000000000000000000000000000" AFTER 12500 ns,
							"000000000000000001000000000" AFTER 12520 ns,
							"000000000000000000000000000" AFTER 12540 ns,
							"000000000000000001000000000" AFTER 12560 ns,
							"000000000000000000000000000" AFTER 12580 ns,
							"000000000000000001000000000" AFTER 12600 ns,
							"000000000000000000000000000" AFTER 12620 ns,
							"000000000000000001000000000" AFTER 12640 ns,
							"000000000000000000000000000" AFTER 12660 ns,
							"000000000000000001000000000" AFTER 12680 ns,
							"000000000000000000000000000" AFTER 12700 ns,
							"000000000000000001000000000" AFTER 12720 ns,
							"000000000000000000000000000" AFTER 12740 ns,
							"000000000000000001000000000" AFTER 12760 ns,
							"000000000000000000000000000" AFTER 12780 ns,
							"000000000000000001000000000" AFTER 12800 ns,
							"000000000000000000000000000" AFTER 12820 ns,
							"000000000000000010000000000" AFTER 12840 ns,
							"000000000000000000000000000" AFTER 12860 ns,
							"000000000000000010000000000" AFTER 12880 ns,
							"000000000000000000000000000" AFTER 12900 ns,
							"000000000000000010000000000" AFTER 12920 ns,
							"000000000000000000000000000" AFTER 12940 ns,
							"000000000000000010000000000" AFTER 12960 ns,
							"000000000000000000000000000" AFTER 12980 ns,
							"000000000000000010000000000" AFTER 13000 ns,
							"000000000000000000000000000" AFTER 13020 ns,
							"000000000000000010000000000" AFTER 13040 ns,
							"000000000000000000000000000" AFTER 13060 ns,
							"000000000000000010000000000" AFTER 13080 ns,
							"000000000000000000000000000" AFTER 13100 ns,
							"000000000000000010000000000" AFTER 13120 ns,
							"000000000000000000000000000" AFTER 13140 ns,
							"000000000000000010000000000" AFTER 13160 ns,
							"000000000000000000000000000" AFTER 13180 ns,
							"000000000000000010000000000" AFTER 13200 ns,
							"000000000000000000000000000" AFTER 13220 ns,
							"000000000000000010000000000" AFTER 13240 ns,
							"000000000000000000000000000" AFTER 13260 ns,
							"000000000000000010000000000" AFTER 13280 ns,
							"000000000000000000000000000" AFTER 13300 ns,
							"000000000000000010000000000" AFTER 13320 ns,
							"000000000000000000000000000" AFTER 13340 ns,
							"000000000000000010000000000" AFTER 13360 ns,
							"000000000000000000000000000" AFTER 13380 ns,
							"000000000000000010000000000" AFTER 13400 ns,
							"000000000000000000000000000" AFTER 13420 ns,
							"000000000000000010000000000" AFTER 13440 ns,
							"000000000000000000000000000" AFTER 13460 ns,
							"000000000000000010000000000" AFTER 13480 ns,
							"000000000000000000000000000" AFTER 13500 ns,
							"000000000000000010000000000" AFTER 13520 ns,
							"000000000000000000000000000" AFTER 13540 ns,
							"000000000000000010000000000" AFTER 13560 ns,
							"000000000000000000000000000" AFTER 13580 ns,
							"000000000000000010000000000" AFTER 13600 ns,
							"000000000000000000000000000" AFTER 13620 ns,
							"000000000000000010000000000" AFTER 13640 ns,
							"000000000000000000000000000" AFTER 13660 ns,
							"000000000000000010000000000" AFTER 13680 ns,
							"000000000000000000000000000" AFTER 13700 ns,
							"000000000000000010000000000" AFTER 13720 ns,
							"000000000000000000000000000" AFTER 13740 ns,
							"000000000000000010000000000" AFTER 13760 ns,
							"000000000000000000000000000" AFTER 13780 ns,
							"000000000000000010000000000" AFTER 13800 ns,
							"000000000000000000000000000" AFTER 13820 ns,
							"000000000000000010000000000" AFTER 13840 ns,
							"000000000000000000000000000" AFTER 13860 ns,
							"000000000000000010000000000" AFTER 13880 ns,
							"000000000000000000000000000" AFTER 13900 ns,
							"000000000000000010000000000" AFTER 13920 ns,
							"000000000000000000000000000" AFTER 13940 ns,
							"000000000000000010000000000" AFTER 13960 ns,
							"000000000000000000000000000" AFTER 13980 ns,
							"000000000000000010000000000" AFTER 14000 ns,
							"000000000000000000000000000" AFTER 14020 ns,
							"000000000000000010000000000" AFTER 14040 ns,
							"000000000000000000000000000" AFTER 14060 ns,
							"000000000000000010000000000" AFTER 14080 ns,
							"000000000000000000000000000" AFTER 14100 ns,
							"000000000000000100000000000" AFTER 14120 ns,
							"000000000000000000000000000" AFTER 14140 ns,
							"000000000000000100000000000" AFTER 14160 ns,
							"000000000000000000000000000" AFTER 14180 ns,
							"000000000000000100000000000" AFTER 14200 ns,
							"000000000000000000000000000" AFTER 14220 ns,
							"000000000000000100000000000" AFTER 14240 ns,
							"000000000000000000000000000" AFTER 14260 ns,
							"000000000000000100000000000" AFTER 14280 ns,
							"000000000000000000000000000" AFTER 14300 ns,
							"000000000000000100000000000" AFTER 14320 ns,
							"000000000000000000000000000" AFTER 14340 ns,
							"000000000000000100000000000" AFTER 14360 ns,
							"000000000000000000000000000" AFTER 14380 ns,
							"000000000000000100000000000" AFTER 14400 ns,
							"000000000000000000000000000" AFTER 14420 ns,
							"000000000000000100000000000" AFTER 14440 ns,
							"000000000000000000000000000" AFTER 14460 ns,
							"000000000000000100000000000" AFTER 14480 ns,
							"000000000000000000000000000" AFTER 14500 ns,
							"000000000000000100000000000" AFTER 14520 ns,
							"000000000000000000000000000" AFTER 14540 ns,
							"000000000000000100000000000" AFTER 14560 ns,
							"000000000000000000000000000" AFTER 14580 ns,
							"000000000000000100000000000" AFTER 14600 ns,
							"000000000000000000000000000" AFTER 14620 ns,
							"000000000000000100000000000" AFTER 14640 ns,
							"000000000000000000000000000" AFTER 14660 ns,
							"000000000000000100000000000" AFTER 14680 ns,
							"000000000000000000000000000" AFTER 14700 ns,
							"000000000000000100000000000" AFTER 14720 ns,
							"000000000000000000000000000" AFTER 14740 ns,
							"000000000000000100000000000" AFTER 14760 ns,
							"000000000000000000000000000" AFTER 14780 ns,
							"000000000000000100000000000" AFTER 14800 ns,
							"000000000000000000000000000" AFTER 14820 ns,
							"000000000000000100000000000" AFTER 14840 ns,
							"000000000000000000000000000" AFTER 14860 ns,
							"000000000000000100000000000" AFTER 14880 ns,
							"000000000000000000000000000" AFTER 14900 ns,
							"000000000000000100000000000" AFTER 14920 ns,
							"000000000000000000000000000" AFTER 14940 ns,
							"000000000000000100000000000" AFTER 14960 ns,
							"000000000000000000000000000" AFTER 14980 ns,
							"000000000000000100000000000" AFTER 15000 ns,
							"000000000000000000000000000" AFTER 15020 ns,
							"000000000000000100000000000" AFTER 15040 ns,
							"000000000000000000000000000" AFTER 15060 ns,
							"000000000000000100000000000" AFTER 15080 ns,
							"000000000000000000000000000" AFTER 15100 ns,
							"000000000000000100000000000" AFTER 15120 ns,
							"000000000000000000000000000" AFTER 15140 ns,
							"000000000000000100000000000" AFTER 15160 ns,
							"000000000000000000000000000" AFTER 15180 ns,
							"000000000000000100000000000" AFTER 15200 ns,
							"000000000000000000000000000" AFTER 15220 ns,
							"000000000000000100000000000" AFTER 15240 ns,
							"000000000000000000000000000" AFTER 15260 ns,
							"000000000000000100000000000" AFTER 15280 ns,
							"000000000000000000000000000" AFTER 15300 ns,
							"000000000000000100000000000" AFTER 15320 ns,
							"000000000000000000000000000" AFTER 15340 ns,
							"000000000000000100000000000" AFTER 15360 ns,
							"000000000000000000000000000" AFTER 15380 ns,
							"000000000000001000000000000" AFTER 15400 ns,
							"000000000000000000000000000" AFTER 15420 ns,
							"000000000000001000000000000" AFTER 15440 ns,
							"000000000000000000000000000" AFTER 15460 ns,
							"000000000000001000000000000" AFTER 15480 ns,
							"000000000000000000000000000" AFTER 15500 ns,
							"000000000000001000000000000" AFTER 15520 ns,
							"000000000000000000000000000" AFTER 15540 ns,
							"000000000000001000000000000" AFTER 15560 ns,
							"000000000000000000000000000" AFTER 15580 ns,
							"000000000000001000000000000" AFTER 15600 ns,
							"000000000000000000000000000" AFTER 15620 ns,
							"000000000000001000000000000" AFTER 15640 ns,
							"000000000000000000000000000" AFTER 15660 ns,
							"000000000000001000000000000" AFTER 15680 ns,
							"000000000000000000000000000" AFTER 15700 ns,
							"000000000000001000000000000" AFTER 15720 ns,
							"000000000000000000000000000" AFTER 15740 ns,
							"000000000000001000000000000" AFTER 15760 ns,
							"000000000000000000000000000" AFTER 15780 ns,
							"000000000000001000000000000" AFTER 15800 ns,
							"000000000000000000000000000" AFTER 15820 ns,
							"000000000000001000000000000" AFTER 15840 ns,
							"000000000000000000000000000" AFTER 15860 ns,
							"000000000000001000000000000" AFTER 15880 ns,
							"000000000000000000000000000" AFTER 15900 ns,
							"000000000000001000000000000" AFTER 15920 ns,
							"000000000000000000000000000" AFTER 15940 ns,
							"000000000000001000000000000" AFTER 15960 ns,
							"000000000000000000000000000" AFTER 15980 ns,
							"000000000000001000000000000" AFTER 16000 ns,
							"000000000000000000000000000" AFTER 16020 ns,
							"000000000000001000000000000" AFTER 16040 ns,
							"000000000000000000000000000" AFTER 16060 ns,
							"000000000000001000000000000" AFTER 16080 ns,
							"000000000000000000000000000" AFTER 16100 ns,
							"000000000000001000000000000" AFTER 16120 ns,
							"000000000000000000000000000" AFTER 16140 ns,
							"000000000000001000000000000" AFTER 16160 ns,
							"000000000000000000000000000" AFTER 16180 ns,
							"000000000000001000000000000" AFTER 16200 ns,
							"000000000000000000000000000" AFTER 16220 ns,
							"000000000000001000000000000" AFTER 16240 ns,
							"000000000000000000000000000" AFTER 16260 ns,
							"000000000000001000000000000" AFTER 16280 ns,
							"000000000000000000000000000" AFTER 16300 ns,
							"000000000000001000000000000" AFTER 16320 ns,
							"000000000000000000000000000" AFTER 16340 ns,
							"000000000000001000000000000" AFTER 16360 ns,
							"000000000000000000000000000" AFTER 16380 ns,
							"000000000000001000000000000" AFTER 16400 ns,
							"000000000000000000000000000" AFTER 16420 ns,
							"000000000000001000000000000" AFTER 16440 ns,
							"000000000000000000000000000" AFTER 16460 ns,
							"000000000000001000000000000" AFTER 16480 ns,
							"000000000000000000000000000" AFTER 16500 ns,
							"000000000000001000000000000" AFTER 16520 ns,
							"000000000000000000000000000" AFTER 16540 ns,
							"000000000000001000000000000" AFTER 16560 ns,
							"000000000000000000000000000" AFTER 16580 ns,
							"000000000000001000000000000" AFTER 16600 ns,
							"000000000000000000000000000" AFTER 16620 ns,
							"000000000000001000000000000" AFTER 16640 ns,
							"000000000000000000000000000" AFTER 16660 ns,
							"000000000000010000000000000" AFTER 16680 ns,
							"000000000000000000000000000" AFTER 16700 ns,
							"000000000000010000000000000" AFTER 16720 ns,
							"000000000000000000000000000" AFTER 16740 ns,
							"000000000000010000000000000" AFTER 16760 ns,
							"000000000000000000000000000" AFTER 16780 ns,
							"000000000000010000000000000" AFTER 16800 ns,
							"000000000000000000000000000" AFTER 16820 ns,
							"000000000000010000000000000" AFTER 16840 ns,
							"000000000000000000000000000" AFTER 16860 ns,
							"000000000000010000000000000" AFTER 16880 ns,
							"000000000000000000000000000" AFTER 16900 ns,
							"000000000000010000000000000" AFTER 16920 ns,
							"000000000000000000000000000" AFTER 16940 ns,
							"000000000000010000000000000" AFTER 16960 ns,
							"000000000000000000000000000" AFTER 16980 ns,
							"000000000000010000000000000" AFTER 17000 ns,
							"000000000000000000000000000" AFTER 17020 ns,
							"000000000000010000000000000" AFTER 17040 ns,
							"000000000000000000000000000" AFTER 17060 ns,
							"000000000000010000000000000" AFTER 17080 ns,
							"000000000000000000000000000" AFTER 17100 ns,
							"000000000000010000000000000" AFTER 17120 ns,
							"000000000000000000000000000" AFTER 17140 ns,
							"000000000000010000000000000" AFTER 17160 ns,
							"000000000000000000000000000" AFTER 17180 ns,
							"000000000000010000000000000" AFTER 17200 ns,
							"000000000000000000000000000" AFTER 17220 ns,
							"000000000000010000000000000" AFTER 17240 ns,
							"000000000000000000000000000" AFTER 17260 ns,
							"000000000000010000000000000" AFTER 17280 ns,
							"000000000000000000000000000" AFTER 17300 ns,
							"000000000000010000000000000" AFTER 17320 ns,
							"000000000000000000000000000" AFTER 17340 ns,
							"000000000000010000000000000" AFTER 17360 ns,
							"000000000000000000000000000" AFTER 17380 ns,
							"000000000000010000000000000" AFTER 17400 ns,
							"000000000000000000000000000" AFTER 17420 ns,
							"000000000000010000000000000" AFTER 17440 ns,
							"000000000000000000000000000" AFTER 17460 ns,
							"000000000000010000000000000" AFTER 17480 ns,
							"000000000000000000000000000" AFTER 17500 ns,
							"000000000000010000000000000" AFTER 17520 ns,
							"000000000000000000000000000" AFTER 17540 ns,
							"000000000000010000000000000" AFTER 17560 ns,
							"000000000000000000000000000" AFTER 17580 ns,
							"000000000000010000000000000" AFTER 17600 ns,
							"000000000000000000000000000" AFTER 17620 ns,
							"000000000000010000000000000" AFTER 17640 ns,
							"000000000000000000000000000" AFTER 17660 ns,
							"000000000000010000000000000" AFTER 17680 ns,
							"000000000000000000000000000" AFTER 17700 ns,
							"000000000000010000000000000" AFTER 17720 ns,
							"000000000000000000000000000" AFTER 17740 ns,
							"000000000000010000000000000" AFTER 17760 ns,
							"000000000000000000000000000" AFTER 17780 ns,
							"000000000000010000000000000" AFTER 17800 ns,
							"000000000000000000000000000" AFTER 17820 ns,
							"000000000000010000000000000" AFTER 17840 ns,
							"000000000000000000000000000" AFTER 17860 ns,
							"000000000000010000000000000" AFTER 17880 ns,
							"000000000000000000000000000" AFTER 17900 ns,
							"000000000000010000000000000" AFTER 17920 ns,
							"000000000000000000000000000" AFTER 17940 ns,
							"000000000000100000000000000" AFTER 17960 ns,
							"000000000000000000000000000" AFTER 17980 ns,
							"000000000000100000000000000" AFTER 18000 ns,
							"000000000000000000000000000" AFTER 18020 ns,
							"000000000000100000000000000" AFTER 18040 ns,
							"000000000000000000000000000" AFTER 18060 ns,
							"000000000000100000000000000" AFTER 18080 ns,
							"000000000000000000000000000" AFTER 18100 ns,
							"000000000000100000000000000" AFTER 18120 ns,
							"000000000000000000000000000" AFTER 18140 ns,
							"000000000000100000000000000" AFTER 18160 ns,
							"000000000000000000000000000" AFTER 18180 ns,
							"000000000000100000000000000" AFTER 18200 ns,
							"000000000000000000000000000" AFTER 18220 ns,
							"000000000000100000000000000" AFTER 18240 ns,
							"000000000000000000000000000" AFTER 18260 ns,
							"000000000000100000000000000" AFTER 18280 ns,
							"000000000000000000000000000" AFTER 18300 ns,
							"000000000000100000000000000" AFTER 18320 ns,
							"000000000000000000000000000" AFTER 18340 ns,
							"000000000000100000000000000" AFTER 18360 ns,
							"000000000000000000000000000" AFTER 18380 ns,
							"000000000000100000000000000" AFTER 18400 ns,
							"000000000000000000000000000" AFTER 18420 ns,
							"000000000000100000000000000" AFTER 18440 ns,
							"000000000000000000000000000" AFTER 18460 ns,
							"000000000000100000000000000" AFTER 18480 ns,
							"000000000000000000000000000" AFTER 18500 ns,
							"000000000000100000000000000" AFTER 18520 ns,
							"000000000000000000000000000" AFTER 18540 ns,
							"000000000000100000000000000" AFTER 18560 ns,
							"000000000000000000000000000" AFTER 18580 ns,
							"000000000000100000000000000" AFTER 18600 ns,
							"000000000000000000000000000" AFTER 18620 ns,
							"000000000000100000000000000" AFTER 18640 ns,
							"000000000000000000000000000" AFTER 18660 ns,
							"000000000000100000000000000" AFTER 18680 ns,
							"000000000000000000000000000" AFTER 18700 ns,
							"000000000000100000000000000" AFTER 18720 ns,
							"000000000000000000000000000" AFTER 18740 ns,
							"000000000000100000000000000" AFTER 18760 ns,
							"000000000000000000000000000" AFTER 18780 ns,
							"000000000000100000000000000" AFTER 18800 ns,
							"000000000000000000000000000" AFTER 18820 ns,
							"000000000000100000000000000" AFTER 18840 ns,
							"000000000000000000000000000" AFTER 18860 ns,
							"000000000000100000000000000" AFTER 18880 ns,
							"000000000000000000000000000" AFTER 18900 ns,
							"000000000000100000000000000" AFTER 18920 ns,
							"000000000000000000000000000" AFTER 18940 ns,
							"000000000000100000000000000" AFTER 18960 ns,
							"000000000000000000000000000" AFTER 18980 ns,
							"000000000000100000000000000" AFTER 19000 ns,
							"000000000000000000000000000" AFTER 19020 ns,
							"000000000000100000000000000" AFTER 19040 ns,
							"000000000000000000000000000" AFTER 19060 ns,
							"000000000000100000000000000" AFTER 19080 ns,
							"000000000000000000000000000" AFTER 19100 ns,
							"000000000000100000000000000" AFTER 19120 ns,
							"000000000000000000000000000" AFTER 19140 ns,
							"000000000000100000000000000" AFTER 19160 ns,
							"000000000000000000000000000" AFTER 19180 ns,
							"000000000000100000000000000" AFTER 19200 ns,
							"000000000000000000000000000" AFTER 19220 ns,
							"000000000001000000000000000" AFTER 19240 ns,
							"000000000000000000000000000" AFTER 19260 ns,
							"000000000001000000000000000" AFTER 19280 ns,
							"000000000000000000000000000" AFTER 19300 ns,
							"000000000001000000000000000" AFTER 19320 ns,
							"000000000000000000000000000" AFTER 19340 ns,
							"000000000001000000000000000" AFTER 19360 ns,
							"000000000000000000000000000" AFTER 19380 ns,
							"000000000001000000000000000" AFTER 19400 ns,
							"000000000000000000000000000" AFTER 19420 ns,
							"000000000001000000000000000" AFTER 19440 ns,
							"000000000000000000000000000" AFTER 19460 ns,
							"000000000001000000000000000" AFTER 19480 ns,
							"000000000000000000000000000" AFTER 19500 ns,
							"000000000001000000000000000" AFTER 19520 ns,
							"000000000000000000000000000" AFTER 19540 ns,
							"000000000001000000000000000" AFTER 19560 ns,
							"000000000000000000000000000" AFTER 19580 ns,
							"000000000001000000000000000" AFTER 19600 ns,
							"000000000000000000000000000" AFTER 19620 ns,
							"000000000001000000000000000" AFTER 19640 ns,
							"000000000000000000000000000" AFTER 19660 ns,
							"000000000001000000000000000" AFTER 19680 ns,
							"000000000000000000000000000" AFTER 19700 ns,
							"000000000001000000000000000" AFTER 19720 ns,
							"000000000000000000000000000" AFTER 19740 ns,
							"000000000001000000000000000" AFTER 19760 ns,
							"000000000000000000000000000" AFTER 19780 ns,
							"000000000001000000000000000" AFTER 19800 ns,
							"000000000000000000000000000" AFTER 19820 ns,
							"000000000001000000000000000" AFTER 19840 ns,
							"000000000000000000000000000" AFTER 19860 ns,
							"000000000001000000000000000" AFTER 19880 ns,
							"000000000000000000000000000" AFTER 19900 ns,
							"000000000001000000000000000" AFTER 19920 ns,
							"000000000000000000000000000" AFTER 19940 ns,
							"000000000001000000000000000" AFTER 19960 ns,
							"000000000000000000000000000" AFTER 19980 ns,
							"000000000001000000000000000" AFTER 20000 ns,
							"000000000000000000000000000" AFTER 20020 ns,
							"000000000001000000000000000" AFTER 20040 ns,
							"000000000000000000000000000" AFTER 20060 ns,
							"000000000001000000000000000" AFTER 20080 ns,
							"000000000000000000000000000" AFTER 20100 ns,
							"000000000001000000000000000" AFTER 20120 ns,
							"000000000000000000000000000" AFTER 20140 ns,
							"000000000001000000000000000" AFTER 20160 ns,
							"000000000000000000000000000" AFTER 20180 ns,
							"000000000001000000000000000" AFTER 20200 ns,
							"000000000000000000000000000" AFTER 20220 ns,
							"000000000001000000000000000" AFTER 20240 ns,
							"000000000000000000000000000" AFTER 20260 ns,
							"000000000001000000000000000" AFTER 20280 ns,
							"000000000000000000000000000" AFTER 20300 ns,
							"000000000001000000000000000" AFTER 20320 ns,
							"000000000000000000000000000" AFTER 20340 ns,
							"000000000001000000000000000" AFTER 20360 ns,
							"000000000000000000000000000" AFTER 20380 ns,
							"000000000001000000000000000" AFTER 20400 ns,
							"000000000000000000000000000" AFTER 20420 ns,
							"000000000001000000000000000" AFTER 20440 ns,
							"000000000000000000000000000" AFTER 20460 ns,
							"000000000001000000000000000" AFTER 20480 ns,
							"000000000000000000000000000" AFTER 20500 ns,
							"000000000010000000000000000" AFTER 20520 ns,
							"000000000000000000000000000" AFTER 20540 ns,
							"000000000010000000000000000" AFTER 20560 ns,
							"000000000000000000000000000" AFTER 20580 ns,
							"000000000010000000000000000" AFTER 20600 ns,
							"000000000000000000000000000" AFTER 20620 ns,
							"000000000010000000000000000" AFTER 20640 ns,
							"000000000000000000000000000" AFTER 20660 ns,
							"000000000010000000000000000" AFTER 20680 ns,
							"000000000000000000000000000" AFTER 20700 ns,
							"000000000010000000000000000" AFTER 20720 ns,
							"000000000000000000000000000" AFTER 20740 ns,
							"000000000010000000000000000" AFTER 20760 ns,
							"000000000000000000000000000" AFTER 20780 ns,
							"000000000010000000000000000" AFTER 20800 ns,
							"000000000000000000000000000" AFTER 20820 ns,
							"000000000010000000000000000" AFTER 20840 ns,
							"000000000000000000000000000" AFTER 20860 ns,
							"000000000010000000000000000" AFTER 20880 ns,
							"000000000000000000000000000" AFTER 20900 ns,
							"000000000010000000000000000" AFTER 20920 ns,
							"000000000000000000000000000" AFTER 20940 ns,
							"000000000010000000000000000" AFTER 20960 ns,
							"000000000000000000000000000" AFTER 20980 ns,
							"000000000010000000000000000" AFTER 21000 ns,
							"000000000000000000000000000" AFTER 21020 ns,
							"000000000010000000000000000" AFTER 21040 ns,
							"000000000000000000000000000" AFTER 21060 ns,
							"000000000010000000000000000" AFTER 21080 ns,
							"000000000000000000000000000" AFTER 21100 ns,
							"000000000010000000000000000" AFTER 21120 ns,
							"000000000000000000000000000" AFTER 21140 ns,
							"000000000010000000000000000" AFTER 21160 ns,
							"000000000000000000000000000" AFTER 21180 ns,
							"000000000010000000000000000" AFTER 21200 ns,
							"000000000000000000000000000" AFTER 21220 ns,
							"000000000010000000000000000" AFTER 21240 ns,
							"000000000000000000000000000" AFTER 21260 ns,
							"000000000010000000000000000" AFTER 21280 ns,
							"000000000000000000000000000" AFTER 21300 ns,
							"000000000010000000000000000" AFTER 21320 ns,
							"000000000000000000000000000" AFTER 21340 ns,
							"000000000010000000000000000" AFTER 21360 ns,
							"000000000000000000000000000" AFTER 21380 ns,
							"000000000010000000000000000" AFTER 21400 ns,
							"000000000000000000000000000" AFTER 21420 ns,
							"000000000010000000000000000" AFTER 21440 ns,
							"000000000000000000000000000" AFTER 21460 ns,
							"000000000010000000000000000" AFTER 21480 ns,
							"000000000000000000000000000" AFTER 21500 ns,
							"000000000010000000000000000" AFTER 21520 ns,
							"000000000000000000000000000" AFTER 21540 ns,
							"000000000010000000000000000" AFTER 21560 ns,
							"000000000000000000000000000" AFTER 21580 ns,
							"000000000010000000000000000" AFTER 21600 ns,
							"000000000000000000000000000" AFTER 21620 ns,
							"000000000010000000000000000" AFTER 21640 ns,
							"000000000000000000000000000" AFTER 21660 ns,
							"000000000010000000000000000" AFTER 21680 ns,
							"000000000000000000000000000" AFTER 21700 ns,
							"000000000010000000000000000" AFTER 21720 ns,
							"000000000000000000000000000" AFTER 21740 ns,
							"000000000010000000000000000" AFTER 21760 ns,
							"000000000000000000000000000" AFTER 21780 ns,
							"000000000100000000000000000" AFTER 21800 ns,
							"000000000000000000000000000" AFTER 21820 ns,
							"000000000100000000000000000" AFTER 21840 ns,
							"000000000000000000000000000" AFTER 21860 ns,
							"000000000100000000000000000" AFTER 21880 ns,
							"000000000000000000000000000" AFTER 21900 ns,
							"000000000100000000000000000" AFTER 21920 ns,
							"000000000000000000000000000" AFTER 21940 ns,
							"000000000100000000000000000" AFTER 21960 ns,
							"000000000000000000000000000" AFTER 21980 ns,
							"000000000100000000000000000" AFTER 22000 ns,
							"000000000000000000000000000" AFTER 22020 ns,
							"000000000100000000000000000" AFTER 22040 ns,
							"000000000000000000000000000" AFTER 22060 ns,
							"000000000100000000000000000" AFTER 22080 ns,
							"000000000000000000000000000" AFTER 22100 ns,
							"000000000100000000000000000" AFTER 22120 ns,
							"000000000000000000000000000" AFTER 22140 ns,
							"000000000100000000000000000" AFTER 22160 ns,
							"000000000000000000000000000" AFTER 22180 ns,
							"000000000100000000000000000" AFTER 22200 ns,
							"000000000000000000000000000" AFTER 22220 ns,
							"000000000100000000000000000" AFTER 22240 ns,
							"000000000000000000000000000" AFTER 22260 ns,
							"000000000100000000000000000" AFTER 22280 ns,
							"000000000000000000000000000" AFTER 22300 ns,
							"000000000100000000000000000" AFTER 22320 ns,
							"000000000000000000000000000" AFTER 22340 ns,
							"000000000100000000000000000" AFTER 22360 ns,
							"000000000000000000000000000" AFTER 22380 ns,
							"000000000100000000000000000" AFTER 22400 ns,
							"000000000000000000000000000" AFTER 22420 ns,
							"000000000100000000000000000" AFTER 22440 ns,
							"000000000000000000000000000" AFTER 22460 ns,
							"000000000100000000000000000" AFTER 22480 ns,
							"000000000000000000000000000" AFTER 22500 ns,
							"000000000100000000000000000" AFTER 22520 ns,
							"000000000000000000000000000" AFTER 22540 ns,
							"000000000100000000000000000" AFTER 22560 ns,
							"000000000000000000000000000" AFTER 22580 ns,
							"000000000100000000000000000" AFTER 22600 ns,
							"000000000000000000000000000" AFTER 22620 ns,
							"000000000100000000000000000" AFTER 22640 ns,
							"000000000000000000000000000" AFTER 22660 ns,
							"000000000100000000000000000" AFTER 22680 ns,
							"000000000000000000000000000" AFTER 22700 ns,
							"000000000100000000000000000" AFTER 22720 ns,
							"000000000000000000000000000" AFTER 22740 ns,
							"000000000100000000000000000" AFTER 22760 ns,
							"000000000000000000000000000" AFTER 22780 ns,
							"000000000100000000000000000" AFTER 22800 ns,
							"000000000000000000000000000" AFTER 22820 ns,
							"000000000100000000000000000" AFTER 22840 ns,
							"000000000000000000000000000" AFTER 22860 ns,
							"000000000100000000000000000" AFTER 22880 ns,
							"000000000000000000000000000" AFTER 22900 ns,
							"000000000100000000000000000" AFTER 22920 ns,
							"000000000000000000000000000" AFTER 22940 ns,
							"000000000100000000000000000" AFTER 22960 ns,
							"000000000000000000000000000" AFTER 22980 ns,
							"000000000100000000000000000" AFTER 23000 ns,
							"000000000000000000000000000" AFTER 23020 ns,
							"000000000100000000000000000" AFTER 23040 ns,
							"000000000000000000000000000" AFTER 23060 ns,
							"000000001000000000000000000" AFTER 23080 ns,
							"000000000000000000000000000" AFTER 23100 ns,
							"000000001000000000000000000" AFTER 23120 ns,
							"000000000000000000000000000" AFTER 23140 ns,
							"000000001000000000000000000" AFTER 23160 ns,
							"000000000000000000000000000" AFTER 23180 ns,
							"000000001000000000000000000" AFTER 23200 ns,
							"000000000000000000000000000" AFTER 23220 ns,
							"000000001000000000000000000" AFTER 23240 ns,
							"000000000000000000000000000" AFTER 23260 ns,
							"000000001000000000000000000" AFTER 23280 ns,
							"000000000000000000000000000" AFTER 23300 ns,
							"000000001000000000000000000" AFTER 23320 ns,
							"000000000000000000000000000" AFTER 23340 ns,
							"000000001000000000000000000" AFTER 23360 ns,
							"000000000000000000000000000" AFTER 23380 ns,
							"000000001000000000000000000" AFTER 23400 ns,
							"000000000000000000000000000" AFTER 23420 ns,
							"000000001000000000000000000" AFTER 23440 ns,
							"000000000000000000000000000" AFTER 23460 ns,
							"000000001000000000000000000" AFTER 23480 ns,
							"000000000000000000000000000" AFTER 23500 ns,
							"000000001000000000000000000" AFTER 23520 ns,
							"000000000000000000000000000" AFTER 23540 ns,
							"000000001000000000000000000" AFTER 23560 ns,
							"000000000000000000000000000" AFTER 23580 ns,
							"000000001000000000000000000" AFTER 23600 ns,
							"000000000000000000000000000" AFTER 23620 ns,
							"000000001000000000000000000" AFTER 23640 ns,
							"000000000000000000000000000" AFTER 23660 ns,
							"000000001000000000000000000" AFTER 23680 ns,
							"000000000000000000000000000" AFTER 23700 ns,
							"000000001000000000000000000" AFTER 23720 ns,
							"000000000000000000000000000" AFTER 23740 ns,
							"000000001000000000000000000" AFTER 23760 ns,
							"000000000000000000000000000" AFTER 23780 ns,
							"000000001000000000000000000" AFTER 23800 ns,
							"000000000000000000000000000" AFTER 23820 ns,
							"000000001000000000000000000" AFTER 23840 ns,
							"000000000000000000000000000" AFTER 23860 ns,
							"000000001000000000000000000" AFTER 23880 ns,
							"000000000000000000000000000" AFTER 23900 ns,
							"000000001000000000000000000" AFTER 23920 ns,
							"000000000000000000000000000" AFTER 23940 ns,
							"000000001000000000000000000" AFTER 23960 ns,
							"000000000000000000000000000" AFTER 23980 ns,
							"000000001000000000000000000" AFTER 24000 ns,
							"000000000000000000000000000" AFTER 24020 ns,
							"000000001000000000000000000" AFTER 24040 ns,
							"000000000000000000000000000" AFTER 24060 ns,
							"000000001000000000000000000" AFTER 24080 ns,
							"000000000000000000000000000" AFTER 24100 ns,
							"000000001000000000000000000" AFTER 24120 ns,
							"000000000000000000000000000" AFTER 24140 ns,
							"000000001000000000000000000" AFTER 24160 ns,
							"000000000000000000000000000" AFTER 24180 ns,
							"000000001000000000000000000" AFTER 24200 ns,
							"000000000000000000000000000" AFTER 24220 ns,
							"000000001000000000000000000" AFTER 24240 ns,
							"000000000000000000000000000" AFTER 24260 ns,
							"000000001000000000000000000" AFTER 24280 ns,
							"000000000000000000000000000" AFTER 24300 ns,
							"000000001000000000000000000" AFTER 24320 ns,
							"000000000000000000000000000" AFTER 24340 ns,
							"000000010000000000000000000" AFTER 24360 ns,
							"000000000000000000000000000" AFTER 24380 ns,
							"000000010000000000000000000" AFTER 24400 ns,
							"000000000000000000000000000" AFTER 24420 ns,
							"000000010000000000000000000" AFTER 24440 ns,
							"000000000000000000000000000" AFTER 24460 ns,
							"000000010000000000000000000" AFTER 24480 ns,
							"000000000000000000000000000" AFTER 24500 ns,
							"000000010000000000000000000" AFTER 24520 ns,
							"000000000000000000000000000" AFTER 24540 ns,
							"000000010000000000000000000" AFTER 24560 ns,
							"000000000000000000000000000" AFTER 24580 ns,
							"000000010000000000000000000" AFTER 24600 ns,
							"000000000000000000000000000" AFTER 24620 ns,
							"000000010000000000000000000" AFTER 24640 ns,
							"000000000000000000000000000" AFTER 24660 ns,
							"000000010000000000000000000" AFTER 24680 ns,
							"000000000000000000000000000" AFTER 24700 ns,
							"000000010000000000000000000" AFTER 24720 ns,
							"000000000000000000000000000" AFTER 24740 ns,
							"000000010000000000000000000" AFTER 24760 ns,
							"000000000000000000000000000" AFTER 24780 ns,
							"000000010000000000000000000" AFTER 24800 ns,
							"000000000000000000000000000" AFTER 24820 ns,
							"000000010000000000000000000" AFTER 24840 ns,
							"000000000000000000000000000" AFTER 24860 ns,
							"000000010000000000000000000" AFTER 24880 ns,
							"000000000000000000000000000" AFTER 24900 ns,
							"000000010000000000000000000" AFTER 24920 ns,
							"000000000000000000000000000" AFTER 24940 ns,
							"000000010000000000000000000" AFTER 24960 ns,
							"000000000000000000000000000" AFTER 24980 ns,
							"000000010000000000000000000" AFTER 25000 ns,
							"000000000000000000000000000" AFTER 25020 ns,
							"000000010000000000000000000" AFTER 25040 ns,
							"000000000000000000000000000" AFTER 25060 ns,
							"000000010000000000000000000" AFTER 25080 ns,
							"000000000000000000000000000" AFTER 25100 ns,
							"000000010000000000000000000" AFTER 25120 ns,
							"000000000000000000000000000" AFTER 25140 ns,
							"000000010000000000000000000" AFTER 25160 ns,
							"000000000000000000000000000" AFTER 25180 ns,
							"000000010000000000000000000" AFTER 25200 ns,
							"000000000000000000000000000" AFTER 25220 ns,
							"000000010000000000000000000" AFTER 25240 ns,
							"000000000000000000000000000" AFTER 25260 ns,
							"000000010000000000000000000" AFTER 25280 ns,
							"000000000000000000000000000" AFTER 25300 ns,
							"000000010000000000000000000" AFTER 25320 ns,
							"000000000000000000000000000" AFTER 25340 ns,
							"000000010000000000000000000" AFTER 25360 ns,
							"000000000000000000000000000" AFTER 25380 ns,
							"000000010000000000000000000" AFTER 25400 ns,
							"000000000000000000000000000" AFTER 25420 ns,
							"000000010000000000000000000" AFTER 25440 ns,
							"000000000000000000000000000" AFTER 25460 ns,
							"000000010000000000000000000" AFTER 25480 ns,
							"000000000000000000000000000" AFTER 25500 ns,
							"000000010000000000000000000" AFTER 25520 ns,
							"000000000000000000000000000" AFTER 25540 ns,
							"000000010000000000000000000" AFTER 25560 ns,
							"000000000000000000000000000" AFTER 25580 ns,
							"000000010000000000000000000" AFTER 25600 ns,
							"000000000000000000000000000" AFTER 25620 ns,
							"000000100000000000000000000" AFTER 25640 ns,
							"000000000000000000000000000" AFTER 25660 ns,
							"000000100000000000000000000" AFTER 25680 ns,
							"000000000000000000000000000" AFTER 25700 ns,
							"000000100000000000000000000" AFTER 25720 ns,
							"000000000000000000000000000" AFTER 25740 ns,
							"000000100000000000000000000" AFTER 25760 ns,
							"000000000000000000000000000" AFTER 25780 ns,
							"000000100000000000000000000" AFTER 25800 ns,
							"000000000000000000000000000" AFTER 25820 ns,
							"000000100000000000000000000" AFTER 25840 ns,
							"000000000000000000000000000" AFTER 25860 ns,
							"000000100000000000000000000" AFTER 25880 ns,
							"000000000000000000000000000" AFTER 25900 ns,
							"000000100000000000000000000" AFTER 25920 ns,
							"000000000000000000000000000" AFTER 25940 ns,
							"000000100000000000000000000" AFTER 25960 ns,
							"000000000000000000000000000" AFTER 25980 ns,
							"000000100000000000000000000" AFTER 26000 ns,
							"000000000000000000000000000" AFTER 26020 ns,
							"000000100000000000000000000" AFTER 26040 ns,
							"000000000000000000000000000" AFTER 26060 ns,
							"000000100000000000000000000" AFTER 26080 ns,
							"000000000000000000000000000" AFTER 26100 ns,
							"000000100000000000000000000" AFTER 26120 ns,
							"000000000000000000000000000" AFTER 26140 ns,
							"000000100000000000000000000" AFTER 26160 ns,
							"000000000000000000000000000" AFTER 26180 ns,
							"000000100000000000000000000" AFTER 26200 ns,
							"000000000000000000000000000" AFTER 26220 ns,
							"000000100000000000000000000" AFTER 26240 ns,
							"000000000000000000000000000" AFTER 26260 ns,
							"000000100000000000000000000" AFTER 26280 ns,
							"000000000000000000000000000" AFTER 26300 ns,
							"000000100000000000000000000" AFTER 26320 ns,
							"000000000000000000000000000" AFTER 26340 ns,
							"000000100000000000000000000" AFTER 26360 ns,
							"000000000000000000000000000" AFTER 26380 ns,
							"000000100000000000000000000" AFTER 26400 ns,
							"000000000000000000000000000" AFTER 26420 ns,
							"000000100000000000000000000" AFTER 26440 ns,
							"000000000000000000000000000" AFTER 26460 ns,
							"000000100000000000000000000" AFTER 26480 ns,
							"000000000000000000000000000" AFTER 26500 ns,
							"000000100000000000000000000" AFTER 26520 ns,
							"000000000000000000000000000" AFTER 26540 ns,
							"000000100000000000000000000" AFTER 26560 ns,
							"000000000000000000000000000" AFTER 26580 ns,
							"000000100000000000000000000" AFTER 26600 ns,
							"000000000000000000000000000" AFTER 26620 ns,
							"000000100000000000000000000" AFTER 26640 ns,
							"000000000000000000000000000" AFTER 26660 ns,
							"000000100000000000000000000" AFTER 26680 ns,
							"000000000000000000000000000" AFTER 26700 ns,
							"000000100000000000000000000" AFTER 26720 ns,
							"000000000000000000000000000" AFTER 26740 ns,
							"000000100000000000000000000" AFTER 26760 ns,
							"000000000000000000000000000" AFTER 26780 ns,
							"000000100000000000000000000" AFTER 26800 ns,
							"000000000000000000000000000" AFTER 26820 ns,
							"000000100000000000000000000" AFTER 26840 ns,
							"000000000000000000000000000" AFTER 26860 ns,
							"000000100000000000000000000" AFTER 26880 ns,
							"000000000000000000000000000" AFTER 26900 ns,
							"000001000000000000000000000" AFTER 26920 ns,
							"000000000000000000000000000" AFTER 26940 ns,
							"000001000000000000000000000" AFTER 26960 ns,
							"000000000000000000000000000" AFTER 26980 ns,
							"000001000000000000000000000" AFTER 27000 ns,
							"000000000000000000000000000" AFTER 27020 ns,
							"000001000000000000000000000" AFTER 27040 ns,
							"000000000000000000000000000" AFTER 27060 ns,
							"000001000000000000000000000" AFTER 27080 ns,
							"000000000000000000000000000" AFTER 27100 ns,
							"000001000000000000000000000" AFTER 27120 ns,
							"000000000000000000000000000" AFTER 27140 ns,
							"000001000000000000000000000" AFTER 27160 ns,
							"000000000000000000000000000" AFTER 27180 ns,
							"000001000000000000000000000" AFTER 27200 ns,
							"000000000000000000000000000" AFTER 27220 ns,
							"000001000000000000000000000" AFTER 27240 ns,
							"000000000000000000000000000" AFTER 27260 ns,
							"000001000000000000000000000" AFTER 27280 ns,
							"000000000000000000000000000" AFTER 27300 ns,
							"000001000000000000000000000" AFTER 27320 ns,
							"000000000000000000000000000" AFTER 27340 ns,
							"000001000000000000000000000" AFTER 27360 ns,
							"000000000000000000000000000" AFTER 27380 ns,
							"000001000000000000000000000" AFTER 27400 ns,
							"000000000000000000000000000" AFTER 27420 ns,
							"000001000000000000000000000" AFTER 27440 ns,
							"000000000000000000000000000" AFTER 27460 ns,
							"000001000000000000000000000" AFTER 27480 ns,
							"000000000000000000000000000" AFTER 27500 ns,
							"000001000000000000000000000" AFTER 27520 ns,
							"000000000000000000000000000" AFTER 27540 ns,
							"000001000000000000000000000" AFTER 27560 ns,
							"000000000000000000000000000" AFTER 27580 ns,
							"000001000000000000000000000" AFTER 27600 ns,
							"000000000000000000000000000" AFTER 27620 ns,
							"000001000000000000000000000" AFTER 27640 ns,
							"000000000000000000000000000" AFTER 27660 ns,
							"000001000000000000000000000" AFTER 27680 ns,
							"000000000000000000000000000" AFTER 27700 ns,
							"000001000000000000000000000" AFTER 27720 ns,
							"000000000000000000000000000" AFTER 27740 ns,
							"000001000000000000000000000" AFTER 27760 ns,
							"000000000000000000000000000" AFTER 27780 ns,
							"000001000000000000000000000" AFTER 27800 ns,
							"000000000000000000000000000" AFTER 27820 ns,
							"000001000000000000000000000" AFTER 27840 ns,
							"000000000000000000000000000" AFTER 27860 ns,
							"000001000000000000000000000" AFTER 27880 ns,
							"000000000000000000000000000" AFTER 27900 ns,
							"000001000000000000000000000" AFTER 27920 ns,
							"000000000000000000000000000" AFTER 27940 ns,
							"000001000000000000000000000" AFTER 27960 ns,
							"000000000000000000000000000" AFTER 27980 ns,
							"000001000000000000000000000" AFTER 28000 ns,
							"000000000000000000000000000" AFTER 28020 ns,
							"000001000000000000000000000" AFTER 28040 ns,
							"000000000000000000000000000" AFTER 28060 ns,
							"000001000000000000000000000" AFTER 28080 ns,
							"000000000000000000000000000" AFTER 28100 ns,
							"000001000000000000000000000" AFTER 28120 ns,
							"000000000000000000000000000" AFTER 28140 ns,
							"000001000000000000000000000" AFTER 28160 ns,
							"000000000000000000000000000" AFTER 28180 ns,
							"000010000000000000000000000" AFTER 28200 ns,
							"000000000000000000000000000" AFTER 28220 ns,
							"000000000000000000000000000" AFTER 28240 ns,
							"000000000000000000000000000" AFTER 28260 ns,
							"000000000000000000000000000" AFTER 28280 ns,
							"000000000000000000000000000" AFTER 28300 ns,
							"000000000000000000000000000" AFTER 28320 ns,
							"000000000000000000000000000" AFTER 28340 ns,
							"000100000000000000000000000" AFTER 28360 ns,
							"000000000000000000000000000" AFTER 28380 ns,
							"000100000000000000000000000" AFTER 28400 ns,
							"000000000000000000000000000" AFTER 28420 ns,
							"000100000000000000000000000" AFTER 28440 ns,
							"000000000000000000000000000" AFTER 28460 ns,
							"000100000000000000000000000" AFTER 28480 ns,
							"000000000000000000000000000" AFTER 28500 ns,
							"000100000000000000000000000" AFTER 28520 ns,
							"000000000000000000000000000" AFTER 28540 ns,
							"000100000000000000000000000" AFTER 28560 ns,
							"000000000000000000000000000" AFTER 28580 ns,
							"000100000000000000000000000" AFTER 28600 ns,
							"000000000000000000000000000" AFTER 28620 ns,
							"000100000000000000000000000" AFTER 28640 ns,
							"000000000000000000000000000" AFTER 28660 ns,
							"000100000000000000000000000" AFTER 28680 ns,
							"000000000000000000000000000" AFTER 28700 ns,
							"000100000000000000000000000" AFTER 28720 ns,
							"000000000000000000000000000" AFTER 28740 ns,
							"000100000000000000000000000" AFTER 28760 ns,
							"000000000000000000000000000" AFTER 28780 ns,
							"000100000000000000000000000" AFTER 28800 ns,
							"000000000000000000000000000" AFTER 28820 ns,
							"000100000000000000000000000" AFTER 28840 ns,
							"000000000000000000000000000" AFTER 28860 ns,
							"000100000000000000000000000" AFTER 28880 ns,
							"000000000000000000000000000" AFTER 28900 ns,
							"000100000000000000000000000" AFTER 28920 ns,
							"000000000000000000000000000" AFTER 28940 ns,
							"000100000000000000000000000" AFTER 28960 ns,
							"000000000000000000000000000" AFTER 28980 ns,
							"000100000000000000000000000" AFTER 29000 ns,
							"000000000000000000000000000" AFTER 29020 ns,
							"000100000000000000000000000" AFTER 29040 ns,
							"000000000000000000000000000" AFTER 29060 ns,
							"000100000000000000000000000" AFTER 29080 ns,
							"000000000000000000000000000" AFTER 29100 ns,
							"000100000000000000000000000" AFTER 29120 ns,
							"000000000000000000000000000" AFTER 29140 ns,
							"000100000000000000000000000" AFTER 29160 ns,
							"000000000000000000000000000" AFTER 29180 ns,
							"000100000000000000000000000" AFTER 29200 ns,
							"000000000000000000000000000" AFTER 29220 ns,
							"000100000000000000000000000" AFTER 29240 ns,
							"000000000000000000000000000" AFTER 29260 ns,
							"000100000000000000000000000" AFTER 29280 ns,
							"000000000000000000000000000" AFTER 29300 ns,
							"000100000000000000000000000" AFTER 29320 ns,
							"000000000000000000000000000" AFTER 29340 ns,
							"000100000000000000000000000" AFTER 29360 ns,
							"000000000000000000000000000" AFTER 29380 ns,
							"000100000000000000000000000" AFTER 29400 ns,
							"000000000000000000000000000" AFTER 29420 ns,
							"000100000000000000000000000" AFTER 29440 ns,
							"000000000000000000000000000" AFTER 29460 ns,
							"000100000000000000000000000" AFTER 29480 ns,
							"000000000000000000000000000" AFTER 29500 ns,
							"000100000000000000000000000" AFTER 29520 ns,
							"000000000000000000000000000" AFTER 29540 ns,
							"000100000000000000000000000" AFTER 29560 ns,
							"000000000000000000000000000" AFTER 29580 ns,
							"000100000000000000000000000" AFTER 29600 ns,
							"000000000000000000000000000" AFTER 29620 ns,
							"001000000000000000000000000" AFTER 29640 ns,
							"000000000000000000000000000" AFTER 29660 ns,
							"100000000000000000000000000" AFTER 29680 ns,
							"000000000000000000000000000" AFTER 29700 ns,
							"100000000000000000000000000" AFTER 29720 ns,
							"000000000000000000000000000" AFTER 29740 ns,
							"100000000000000000000000000" AFTER 29760 ns,
							"000000000000000000000000000" AFTER 29780 ns,
							"100000000000000000000000000" AFTER 29800 ns,
							"000000000000000000000000000" AFTER 29820 ns,
							"100000000000000000000000000" AFTER 29840 ns,
							"000000000000000000000000000" AFTER 29860 ns,
							"100000000000000000000000000" AFTER 29880 ns,
							"000000000000000000000000000" AFTER 29900 ns,
							"100000000000000000000000000" AFTER 29920 ns,
							"000000000000000000000000000" AFTER 29940 ns,
							"100000000000000000000000000" AFTER 29960 ns,
							"000000000000000000000000000" AFTER 29980 ns,
							"100000000000000000000000000" AFTER 30000 ns,
							"000000000000000000000000000" AFTER 30020 ns,
							"100000000000000000000000000" AFTER 30040 ns,
							"000000000000000000000000000" AFTER 30060 ns,
							"100000000000000000000000000" AFTER 30080 ns,
							"000000000000000000000000000" AFTER 30100 ns,
							"100000000000000000000000000" AFTER 30120 ns,
							"000000000000000000000000000" AFTER 30140 ns,
							"100000000000000000000000000" AFTER 30160 ns,
							"000000000000000000000000000" AFTER 30180 ns,
							"100000000000000000000000000" AFTER 30200 ns,
							"000000000000000000000000000" AFTER 30220 ns,
							"100000000000000000000000000" AFTER 30240 ns,
							"000000000000000000000000000" AFTER 30260 ns,
							"100000000000000000000000000" AFTER 30280 ns,
							"000000000000000000000000000" AFTER 30300 ns,
							"100000000000000000000000000" AFTER 30320 ns,
							"000000000000000000000000000" AFTER 30340 ns,
							"100000000000000000000000000" AFTER 30360 ns,
							"000000000000000000000000000" AFTER 30380 ns,
							"100000000000000000000000000" AFTER 30400 ns,
							"000000000000000000000000000" AFTER 30420 ns,
							"100000000000000000000000000" AFTER 30440 ns,
							"000000000000000000000000000" AFTER 30460 ns,
							"100000000000000000000000000" AFTER 30480 ns,
							"000000000000000000000000000" AFTER 30500 ns,
							"100000000000000000000000000" AFTER 30520 ns,
							"000000000000000000000000000" AFTER 30540 ns,
							"100000000000000000000000000" AFTER 30560 ns,
							"000000000000000000000000000" AFTER 30580 ns,
							"100000000000000000000000000" AFTER 30600 ns,
							"000000000000000000000000000" AFTER 30620 ns,
							"100000000000000000000000000" AFTER 30640 ns,
							"000000000000000000000000000" AFTER 30660 ns,
							"100000000000000000000000000" AFTER 30680 ns,
							"000000000000000000000000000" AFTER 30700 ns,
							"100000000000000000000000000" AFTER 30720 ns,
							"000000000000000000000000000" AFTER 30740 ns,
							"100000000000000000000000000" AFTER 30760 ns,
							"000000000000000000000000000" AFTER 30780 ns,
							"100000000000000000000000000" AFTER 30800 ns,
							"000000000000000000000000000" AFTER 30820 ns,
							"100000000000000000000000000" AFTER 30840 ns,
							"000000000000000000000000000" AFTER 30860 ns,
							"100000000000000000000000000" AFTER 30880 ns,
							"000000000000000000000000000" AFTER 30900 ns,
							"100000000000000000000000000" AFTER 30920 ns,
							"000000000000000000000000000" AFTER 30940 ns,
							"010000000000000000000000000" AFTER 30960 ns;

IrRegisters <= "00000000000000000000000000000000" AFTER 00020 ns,
					"00000000000000000000000000000000" AFTER 00040 ns,
					"00000000000000000000000000000000" AFTER 00060 ns,
					"00000000000000000000000010000000" AFTER 00080 ns,
					"00000000000000000000000000000000" AFTER 00100 ns,
					"00000000000000000000000100000000" AFTER 00120 ns,
					"00000000000000000000000000000000" AFTER 00140 ns,
					"00000000000000000000000110000000" AFTER 00160 ns,
					"00000000000000000000000000000000" AFTER 00180 ns,
					"00000000000000000000001000000000" AFTER 00200 ns,
					"00000000000000000000000000000000" AFTER 00220 ns,
					"00000000000000000000001010000000" AFTER 00240 ns,
					"00000000000000000000000000000000" AFTER 00260 ns,
					"00000000000000000000001100000000" AFTER 00280 ns,
					"00000000000000000000000000000000" AFTER 00300 ns,
					"00000000000000000000001110000000" AFTER 00320 ns,
					"00000000000000000000000000000000" AFTER 00340 ns,
					"00000000000000000000010000000000" AFTER 00360 ns,
					"00000000000000000000000000000000" AFTER 00380 ns,
					"00000000000000000000010010000000" AFTER 00400 ns,
					"00000000000000000000000000000000" AFTER 00420 ns,
					"00000000000000000000010100000000" AFTER 00440 ns,
					"00000000000000000000000000000000" AFTER 00460 ns,
					"00000000000000000000010110000000" AFTER 00480 ns,
					"00000000000000000000000000000000" AFTER 00500 ns,
					"00000000000000000000011000000000" AFTER 00520 ns,
					"00000000000000000000000000000000" AFTER 00540 ns,
					"00000000000000000000011010000000" AFTER 00560 ns,
					"00000000000000000000000000000000" AFTER 00580 ns,
					"00000000000000000000011100000000" AFTER 00600 ns,
					"00000000000000000000000000000000" AFTER 00620 ns,
					"00000000000000000000011110000000" AFTER 00640 ns,
					"00000000000000000000000000000000" AFTER 00660 ns,
					"00000000000000000000100000000000" AFTER 00680 ns,
					"00000000000000000000000000000000" AFTER 00700 ns,
					"00000000000000000000100010000000" AFTER 00720 ns,
					"00000000000000000000000000000000" AFTER 00740 ns,
					"00000000000000000000100100000000" AFTER 00760 ns,
					"00000000000000000000000000000000" AFTER 00780 ns,
					"00000000000000000000100110000000" AFTER 00800 ns,
					"00000000000000000000000000000000" AFTER 00820 ns,
					"00000000000000000000101000000000" AFTER 00840 ns,
					"00000000000000000000000000000000" AFTER 00860 ns,
					"00000000000000000000101010000000" AFTER 00880 ns,
					"00000000000000000000000000000000" AFTER 00900 ns,
					"00000000000000000000101100000000" AFTER 00920 ns,
					"00000000000000000000000000000000" AFTER 00940 ns,
					"00000000000000000000101110000000" AFTER 00960 ns,
					"00000000000000000000000000000000" AFTER 00980 ns,
					"00000000000000000000110000000000" AFTER 01000 ns,
					"00000000000000000000000000000000" AFTER 01020 ns,
					"00000000000000000000110010000000" AFTER 01040 ns,
					"00000000000000000000000000000000" AFTER 01060 ns,
					"00000000000000000000110100000000" AFTER 01080 ns,
					"00000000000000000000000000000000" AFTER 01100 ns,
					"00000000000000000000110110000000" AFTER 01120 ns,
					"00000000000000000000000000000000" AFTER 01140 ns,
					"00000000000000000000111000000000" AFTER 01160 ns,
					"00000000000000000000000000000000" AFTER 01180 ns,
					"00000000000000000000111010000000" AFTER 01200 ns,
					"00000000000000000000000000000000" AFTER 01220 ns,
					"00000000000000000000111100000000" AFTER 01240 ns,
					"00000000000000000000000000000000" AFTER 01260 ns,
					"00000000000000000000111110000000" AFTER 01280 ns,
					"00000000000000000000000000000000" AFTER 01300 ns,
					"00000000010010110100000000000000" AFTER 01320 ns,
					"00000000000000000000000000000000" AFTER 01340 ns,
					"00000000010010101111000010000000" AFTER 01360 ns,
					"00000000000000000000000000000000" AFTER 01380 ns,
					"00000000010010101010000100000000" AFTER 01400 ns,
					"00000000000000000000000000000000" AFTER 01420 ns,
					"00000000010010100101000110000000" AFTER 01440 ns,
					"00000000000000000000000000000000" AFTER 01460 ns,
					"00000000010010100010001000000000" AFTER 01480 ns,
					"00000000000000000000000000000000" AFTER 01500 ns,
					"00000000010001011111001010000000" AFTER 01520 ns,
					"00000000000000000000000000000000" AFTER 01540 ns,
					"00000000010001011100001100000000" AFTER 01560 ns,
					"00000000000000000000000000000000" AFTER 01580 ns,
					"00000000010001010111001110000000" AFTER 01600 ns,
					"00000000000000000000000000000000" AFTER 01620 ns,
					"00000000010001010010010000000000" AFTER 01640 ns,
					"00000000000000000000000000000000" AFTER 01660 ns,
					"00000000010010001101010010000000" AFTER 01680 ns,
					"00000000000000000000000000000000" AFTER 01700 ns,
					"00000000010010001010010100000000" AFTER 01720 ns,
					"00000000000000000000000000000000" AFTER 01740 ns,
					"00000000010010000111010110000000" AFTER 01760 ns,
					"00000000000000000000000000000000" AFTER 01780 ns,
					"00000000010010000100011000000000" AFTER 01800 ns,
					"00000000000000000000000000000000" AFTER 01820 ns,
					"00000000010001111111011010000000" AFTER 01840 ns,
					"00000000000000000000000000000000" AFTER 01860 ns,
					"00000000010001111010011100000000" AFTER 01880 ns,
					"00000000000000000000000000000000" AFTER 01900 ns,
					"00000000010001110101011110000000" AFTER 01920 ns,
					"00000000000000000000000000000000" AFTER 01940 ns,
					"00000000010001110010100000000000" AFTER 01960 ns,
					"00000000000000000000000000000000" AFTER 01980 ns,
					"00000000010001101111100010000000" AFTER 02000 ns,
					"00000000000000000000000000000000" AFTER 02020 ns,
					"00000000010001101100100100000000" AFTER 02040 ns,
					"00000000000000000000000000000000" AFTER 02060 ns,
					"00000000010001100111100110000000" AFTER 02080 ns,
					"00000000000000000000000000000000" AFTER 02100 ns,
					"00000000010001100010101000000000" AFTER 02120 ns,
					"00000000000000000000000000000000" AFTER 02140 ns,
					"00000000010001011101101010000000" AFTER 02160 ns,
					"00000000000000000000000000000000" AFTER 02180 ns,
					"00000000010001011010101100000000" AFTER 02200 ns,
					"00000000000000000000000000000000" AFTER 02220 ns,
					"00000000010001010111101110000000" AFTER 02240 ns,
					"00000000000000000000000000000000" AFTER 02260 ns,
					"00000000010001010100110000000000" AFTER 02280 ns,
					"00000000000000000000000000000000" AFTER 02300 ns,
					"00000000010001001111110010000000" AFTER 02320 ns,
					"00000000000000000000000000000000" AFTER 02340 ns,
					"00000000010001001010110100000000" AFTER 02360 ns,
					"00000000000000000000000000000000" AFTER 02380 ns,
					"00000000010001000101110110000000" AFTER 02400 ns,
					"00000000000000000000000000000000" AFTER 02420 ns,
					"00000000010001000010111000000000" AFTER 02440 ns,
					"00000000000000000000000000000000" AFTER 02460 ns,
					"00000000010000111111111010000000" AFTER 02480 ns,
					"00000000000000000000000000000000" AFTER 02500 ns,
					"00000000010000111100111100000000" AFTER 02520 ns,
					"00000000000000000000000000000000" AFTER 02540 ns,
					"00000000010000110111111110000000" AFTER 02560 ns,
					"00000000000000000000000000000000" AFTER 02580 ns,
					"00000000000000000000000000000000" AFTER 02600 ns,
					"00000000000000000000000000000000" AFTER 02620 ns,
					"00000000000000001000000000000000" AFTER 02640 ns,
					"00000000000000000000000000000000" AFTER 02660 ns,
					"00000000000000010000000000000000" AFTER 02680 ns,
					"00000000000000000000000000000000" AFTER 02700 ns,
					"00000000000000011000000000000000" AFTER 02720 ns,
					"00000000000000000000000000000000" AFTER 02740 ns,
					"00000000000000100000000000000000" AFTER 02760 ns,
					"00000000000000000000000000000000" AFTER 02780 ns,
					"00000000000000101000000000000000" AFTER 02800 ns,
					"00000000000000000000000000000000" AFTER 02820 ns,
					"00000000000000110000000000000000" AFTER 02840 ns,
					"00000000000000000000000000000000" AFTER 02860 ns,
					"00000000000000111000000000000000" AFTER 02880 ns,
					"00000000000000000000000000000000" AFTER 02900 ns,
					"00000000000001000000000000000000" AFTER 02920 ns,
					"00000000000000000000000000000000" AFTER 02940 ns,
					"00000000000001001000000000000000" AFTER 02960 ns,
					"00000000000000000000000000000000" AFTER 02980 ns,
					"00000000000001010000000000000000" AFTER 03000 ns,
					"00000000000000000000000000000000" AFTER 03020 ns,
					"00000000000001011000000000000000" AFTER 03040 ns,
					"00000000000000000000000000000000" AFTER 03060 ns,
					"00000000000001100000000000000000" AFTER 03080 ns,
					"00000000000000000000000000000000" AFTER 03100 ns,
					"00000000000001101000000000000000" AFTER 03120 ns,
					"00000000000000000000000000000000" AFTER 03140 ns,
					"00000000000001110000000000000000" AFTER 03160 ns,
					"00000000000000000000000000000000" AFTER 03180 ns,
					"00000000000001111000000000000000" AFTER 03200 ns,
					"00000000000000000000000000000000" AFTER 03220 ns,
					"00000000000010000000000000000000" AFTER 03240 ns,
					"00000000000000000000000000000000" AFTER 03260 ns,
					"00000000000010001000000000000000" AFTER 03280 ns,
					"00000000000000000000000000000000" AFTER 03300 ns,
					"00000000000010010000000000000000" AFTER 03320 ns,
					"00000000000000000000000000000000" AFTER 03340 ns,
					"00000000000010011000000000000000" AFTER 03360 ns,
					"00000000000000000000000000000000" AFTER 03380 ns,
					"00000000000010100000000000000000" AFTER 03400 ns,
					"00000000000000000000000000000000" AFTER 03420 ns,
					"00000000000010101000000000000000" AFTER 03440 ns,
					"00000000000000000000000000000000" AFTER 03460 ns,
					"00000000000010110000000000000000" AFTER 03480 ns,
					"00000000000000000000000000000000" AFTER 03500 ns,
					"00000000000010111000000000000000" AFTER 03520 ns,
					"00000000000000000000000000000000" AFTER 03540 ns,
					"00000000000011000000000000000000" AFTER 03560 ns,
					"00000000000000000000000000000000" AFTER 03580 ns,
					"00000000000011001000000000000000" AFTER 03600 ns,
					"00000000000000000000000000000000" AFTER 03620 ns,
					"00000000000011010000000000000000" AFTER 03640 ns,
					"00000000000000000000000000000000" AFTER 03660 ns,
					"00000000000011011000000000000000" AFTER 03680 ns,
					"00000000000000000000000000000000" AFTER 03700 ns,
					"00000000000011100000000000000000" AFTER 03720 ns,
					"00000000000000000000000000000000" AFTER 03740 ns,
					"00000000000011101000000000000000" AFTER 03760 ns,
					"00000000000000000000000000000000" AFTER 03780 ns,
					"00000000000011110000000000000000" AFTER 03800 ns,
					"00000000000000000000000000000000" AFTER 03820 ns,
					"00000000000011111000000000000000" AFTER 03840 ns,
					"00000000000000000000000000000000" AFTER 03860 ns,
					"00000001111100000000000000000000" AFTER 03880 ns,
					"00000000000000000000000000000000" AFTER 03900 ns,
					"00000001111000001000000000000000" AFTER 03920 ns,
					"00000000000000000000000000000000" AFTER 03940 ns,
					"00000001110100010000000000000000" AFTER 03960 ns,
					"00000000000000000000000000000000" AFTER 03980 ns,
					"00000001110000011000000000000000" AFTER 04000 ns,
					"00000000000000000000000000000000" AFTER 04020 ns,
					"00000001101100100000000000000000" AFTER 04040 ns,
					"00000000000000000000000000000000" AFTER 04060 ns,
					"00000001101000101000000000000000" AFTER 04080 ns,
					"00000000000000000000000000000000" AFTER 04100 ns,
					"00000001100100110000000000000000" AFTER 04120 ns,
					"00000000000000000000000000000000" AFTER 04140 ns,
					"00000001100000111000000000000000" AFTER 04160 ns,
					"00000000000000000000000000000000" AFTER 04180 ns,
					"00000001011101000000000000000000" AFTER 04200 ns,
					"00000000000000000000000000000000" AFTER 04220 ns,
					"00000001011001001000000000000000" AFTER 04240 ns,
					"00000000000000000000000000000000" AFTER 04260 ns,
					"00000001010101010000000000000000" AFTER 04280 ns,
					"00000000000000000000000000000000" AFTER 04300 ns,
					"00000001010001011000000000000000" AFTER 04320 ns,
					"00000000000000000000000000000000" AFTER 04340 ns,
					"00000001001101100000000000000000" AFTER 04360 ns,
					"00000000000000000000000000000000" AFTER 04380 ns,
					"00000001001001101000000000000000" AFTER 04400 ns,
					"00000000000000000000000000000000" AFTER 04420 ns,
					"00000001000101110000000000000000" AFTER 04440 ns,
					"00000000000000000000000000000000" AFTER 04460 ns,
					"00000001000001111000000000000000" AFTER 04480 ns,
					"00000000000000000000000000000000" AFTER 04500 ns,
					"00000000111110000000000000000000" AFTER 04520 ns,
					"00000000000000000000000000000000" AFTER 04540 ns,
					"00000000111010001000000000000000" AFTER 04560 ns,
					"00000000000000000000000000000000" AFTER 04580 ns,
					"00000000110110010000000000000000" AFTER 04600 ns,
					"00000000000000000000000000000000" AFTER 04620 ns,
					"00000000110010011000000000000000" AFTER 04640 ns,
					"00000000000000000000000000000000" AFTER 04660 ns,
					"00000000101110100000000000000000" AFTER 04680 ns,
					"00000000000000000000000000000000" AFTER 04700 ns,
					"00000000101010101000000000000000" AFTER 04720 ns,
					"00000000000000000000000000000000" AFTER 04740 ns,
					"00000000100110110000000000000000" AFTER 04760 ns,
					"00000000000000000000000000000000" AFTER 04780 ns,
					"00000000100010111000000000000000" AFTER 04800 ns,
					"00000000000000000000000000000000" AFTER 04820 ns,
					"00000000011111000000000000000000" AFTER 04840 ns,
					"00000000000000000000000000000000" AFTER 04860 ns,
					"00000000011011001000000000000000" AFTER 04880 ns,
					"00000000000000000000000000000000" AFTER 04900 ns,
					"00000000010111010000000000000000" AFTER 04920 ns,
					"00000000000000000000000000000000" AFTER 04940 ns,
					"00000000010011011000000000000000" AFTER 04960 ns,
					"00000000000000000000000000000000" AFTER 04980 ns,
					"00000000001111100000000000000000" AFTER 05000 ns,
					"00000000000000000000000000000000" AFTER 05020 ns,
					"00000000001011101000000000000000" AFTER 05040 ns,
					"00000000000000000000000000000000" AFTER 05060 ns,
					"00000000000111110000000000000000" AFTER 05080 ns,
					"00000000000000000000000000000000" AFTER 05100 ns,
					"00000000000011111000000000000000" AFTER 05120 ns,
					"00000000000000000000000000000000" AFTER 05140 ns,
					"00000000000000000000000000000000" AFTER 05160 ns,
					"00000000000000000000000000000000" AFTER 05180 ns,
					"00000000000000000000000010000000" AFTER 05200 ns,
					"00000000000000000000000000000000" AFTER 05220 ns,
					"00000000000000000000000100000000" AFTER 05240 ns,
					"00000000000000000000000000000000" AFTER 05260 ns,
					"00000000000000000000000110000000" AFTER 05280 ns,
					"00000000000000000000000000000000" AFTER 05300 ns,
					"00000000000000000000001000000000" AFTER 05320 ns,
					"00000000000000000000000000000000" AFTER 05340 ns,
					"00000000000000000000001010000000" AFTER 05360 ns,
					"00000000000000000000000000000000" AFTER 05380 ns,
					"00000000000000000000001100000000" AFTER 05400 ns,
					"00000000000000000000000000000000" AFTER 05420 ns,
					"00000000000000000000001110000000" AFTER 05440 ns,
					"00000000000000000000000000000000" AFTER 05460 ns,
					"00000000000000000000010000000000" AFTER 05480 ns,
					"00000000000000000000000000000000" AFTER 05500 ns,
					"00000000000000000000010010000000" AFTER 05520 ns,
					"00000000000000000000000000000000" AFTER 05540 ns,
					"00000000000000000000010100000000" AFTER 05560 ns,
					"00000000000000000000000000000000" AFTER 05580 ns,
					"00000000000000000000010110000000" AFTER 05600 ns,
					"00000000000000000000000000000000" AFTER 05620 ns,
					"00000000000000000000011000000000" AFTER 05640 ns,
					"00000000000000000000000000000000" AFTER 05660 ns,
					"00000000000000000000011010000000" AFTER 05680 ns,
					"00000000000000000000000000000000" AFTER 05700 ns,
					"00000000000000000000011100000000" AFTER 05720 ns,
					"00000000000000000000000000000000" AFTER 05740 ns,
					"00000000000000000000011110000000" AFTER 05760 ns,
					"00000000000000000000000000000000" AFTER 05780 ns,
					"00000000000000000000100000000000" AFTER 05800 ns,
					"00000000000000000000000000000000" AFTER 05820 ns,
					"00000000000000000000100010000000" AFTER 05840 ns,
					"00000000000000000000000000000000" AFTER 05860 ns,
					"00000000000000000000100100000000" AFTER 05880 ns,
					"00000000000000000000000000000000" AFTER 05900 ns,
					"00000000000000000000100110000000" AFTER 05920 ns,
					"00000000000000000000000000000000" AFTER 05940 ns,
					"00000000000000000000101000000000" AFTER 05960 ns,
					"00000000000000000000000000000000" AFTER 05980 ns,
					"00000000000000000000101010000000" AFTER 06000 ns,
					"00000000000000000000000000000000" AFTER 06020 ns,
					"00000000000000000000101100000000" AFTER 06040 ns,
					"00000000000000000000000000000000" AFTER 06060 ns,
					"00000000000000000000101110000000" AFTER 06080 ns,
					"00000000000000000000000000000000" AFTER 06100 ns,
					"00000000000000000000110000000000" AFTER 06120 ns,
					"00000000000000000000000000000000" AFTER 06140 ns,
					"00000000000000000000110010000000" AFTER 06160 ns,
					"00000000000000000000000000000000" AFTER 06180 ns,
					"00000000000000000000110100000000" AFTER 06200 ns,
					"00000000000000000000000000000000" AFTER 06220 ns,
					"00000000000000000000110110000000" AFTER 06240 ns,
					"00000000000000000000000000000000" AFTER 06260 ns,
					"00000000000000000000111000000000" AFTER 06280 ns,
					"00000000000000000000000000000000" AFTER 06300 ns,
					"00000000000000000000111010000000" AFTER 06320 ns,
					"00000000000000000000000000000000" AFTER 06340 ns,
					"00000000000000000000111100000000" AFTER 06360 ns,
					"00000000000000000000000000000000" AFTER 06380 ns,
					"00000000000000000000111110000000" AFTER 06400 ns,
					"00000000000000000000000000000000" AFTER 06420 ns,
					"00000001111100000000000000000000" AFTER 06440 ns,
					"00000000000000000000000000000000" AFTER 06460 ns,
					"00000001111000001000000000000000" AFTER 06480 ns,
					"00000000000000000000000000000000" AFTER 06500 ns,
					"00000001110100010000000000000000" AFTER 06520 ns,
					"00000000000000000000000000000000" AFTER 06540 ns,
					"00000001110000011000000000000000" AFTER 06560 ns,
					"00000000000000000000000000000000" AFTER 06580 ns,
					"00000001101100100000000000000000" AFTER 06600 ns,
					"00000000000000000000000000000000" AFTER 06620 ns,
					"00000001101000101000000000000000" AFTER 06640 ns,
					"00000000000000000000000000000000" AFTER 06660 ns,
					"00000001100100110000000000000000" AFTER 06680 ns,
					"00000000000000000000000000000000" AFTER 06700 ns,
					"00000001100000111000000000000000" AFTER 06720 ns,
					"00000000000000000000000000000000" AFTER 06740 ns,
					"00000001011101000000000000000000" AFTER 06760 ns,
					"00000000000000000000000000000000" AFTER 06780 ns,
					"00000001011001001000000000000000" AFTER 06800 ns,
					"00000000000000000000000000000000" AFTER 06820 ns,
					"00000001010101010000000000000000" AFTER 06840 ns,
					"00000000000000000000000000000000" AFTER 06860 ns,
					"00000001010001011000000000000000" AFTER 06880 ns,
					"00000000000000000000000000000000" AFTER 06900 ns,
					"00000001001101100000000000000000" AFTER 06920 ns,
					"00000000000000000000000000000000" AFTER 06940 ns,
					"00000001001001101000000000000000" AFTER 06960 ns,
					"00000000000000000000000000000000" AFTER 06980 ns,
					"00000001000101110000000000000000" AFTER 07000 ns,
					"00000000000000000000000000000000" AFTER 07020 ns,
					"00000001000001111000000000000000" AFTER 07040 ns,
					"00000000000000000000000000000000" AFTER 07060 ns,
					"00000000111110000000000000000000" AFTER 07080 ns,
					"00000000000000000000000000000000" AFTER 07100 ns,
					"00000000111010001000000000000000" AFTER 07120 ns,
					"00000000000000000000000000000000" AFTER 07140 ns,
					"00000000110110010000000000000000" AFTER 07160 ns,
					"00000000000000000000000000000000" AFTER 07180 ns,
					"00000000110010011000000000000000" AFTER 07200 ns,
					"00000000000000000000000000000000" AFTER 07220 ns,
					"00000000101110100000000000000000" AFTER 07240 ns,
					"00000000000000000000000000000000" AFTER 07260 ns,
					"00000000101010101000000000000000" AFTER 07280 ns,
					"00000000000000000000000000000000" AFTER 07300 ns,
					"00000000100110110000000000000000" AFTER 07320 ns,
					"00000000000000000000000000000000" AFTER 07340 ns,
					"00000000100010111000000000000000" AFTER 07360 ns,
					"00000000000000000000000000000000" AFTER 07380 ns,
					"00000000011111000000000000000000" AFTER 07400 ns,
					"00000000000000000000000000000000" AFTER 07420 ns,
					"00000000011011001000000000000000" AFTER 07440 ns,
					"00000000000000000000000000000000" AFTER 07460 ns,
					"00000000010111010000000000000000" AFTER 07480 ns,
					"00000000000000000000000000000000" AFTER 07500 ns,
					"00000000010011011000000000000000" AFTER 07520 ns,
					"00000000000000000000000000000000" AFTER 07540 ns,
					"00000000001111100000000000000000" AFTER 07560 ns,
					"00000000000000000000000000000000" AFTER 07580 ns,
					"00000000001011101000000000000000" AFTER 07600 ns,
					"00000000000000000000000000000000" AFTER 07620 ns,
					"00000000000111110000000000000000" AFTER 07640 ns,
					"00000000000000000000000000000000" AFTER 07660 ns,
					"00000000000011111000000000000000" AFTER 07680 ns,
					"00000000000000000000000000000000" AFTER 07700 ns,
					"00000000000000000000000000000000" AFTER 07720 ns,
					"00000000000000000000000000000000" AFTER 07740 ns,
					"00000000000000000000000010000000" AFTER 07760 ns,
					"00000000000000000000000000000000" AFTER 07780 ns,
					"00000000000000000000000100000000" AFTER 07800 ns,
					"00000000000000000000000000000000" AFTER 07820 ns,
					"00000000000000000000000110000000" AFTER 07840 ns,
					"00000000000000000000000000000000" AFTER 07860 ns,
					"00000000000000000000001000000000" AFTER 07880 ns,
					"00000000000000000000000000000000" AFTER 07900 ns,
					"00000000000000000000001010000000" AFTER 07920 ns,
					"00000000000000000000000000000000" AFTER 07940 ns,
					"00000000000000000000001100000000" AFTER 07960 ns,
					"00000000000000000000000000000000" AFTER 07980 ns,
					"00000000000000000000001110000000" AFTER 08000 ns,
					"00000000000000000000000000000000" AFTER 08020 ns,
					"00000000000000000000010000000000" AFTER 08040 ns,
					"00000000000000000000000000000000" AFTER 08060 ns,
					"00000000000000000000010010000000" AFTER 08080 ns,
					"00000000000000000000000000000000" AFTER 08100 ns,
					"00000000000000000000010100000000" AFTER 08120 ns,
					"00000000000000000000000000000000" AFTER 08140 ns,
					"00000000000000000000010110000000" AFTER 08160 ns,
					"00000000000000000000000000000000" AFTER 08180 ns,
					"00000000000000000000011000000000" AFTER 08200 ns,
					"00000000000000000000000000000000" AFTER 08220 ns,
					"00000000000000000000011010000000" AFTER 08240 ns,
					"00000000000000000000000000000000" AFTER 08260 ns,
					"00000000000000000000011100000000" AFTER 08280 ns,
					"00000000000000000000000000000000" AFTER 08300 ns,
					"00000000000000000000011110000000" AFTER 08320 ns,
					"00000000000000000000000000000000" AFTER 08340 ns,
					"00000000000000000000100000000000" AFTER 08360 ns,
					"00000000000000000000000000000000" AFTER 08380 ns,
					"00000000000000000000100010000000" AFTER 08400 ns,
					"00000000000000000000000000000000" AFTER 08420 ns,
					"00000000000000000000100100000000" AFTER 08440 ns,
					"00000000000000000000000000000000" AFTER 08460 ns,
					"00000000000000000000100110000000" AFTER 08480 ns,
					"00000000000000000000000000000000" AFTER 08500 ns,
					"00000000000000000000101000000000" AFTER 08520 ns,
					"00000000000000000000000000000000" AFTER 08540 ns,
					"00000000000000000000101010000000" AFTER 08560 ns,
					"00000000000000000000000000000000" AFTER 08580 ns,
					"00000000000000000000101100000000" AFTER 08600 ns,
					"00000000000000000000000000000000" AFTER 08620 ns,
					"00000000000000000000101110000000" AFTER 08640 ns,
					"00000000000000000000000000000000" AFTER 08660 ns,
					"00000000000000000000110000000000" AFTER 08680 ns,
					"00000000000000000000000000000000" AFTER 08700 ns,
					"00000000000000000000110010000000" AFTER 08720 ns,
					"00000000000000000000000000000000" AFTER 08740 ns,
					"00000000000000000000110100000000" AFTER 08760 ns,
					"00000000000000000000000000000000" AFTER 08780 ns,
					"00000000000000000000110110000000" AFTER 08800 ns,
					"00000000000000000000000000000000" AFTER 08820 ns,
					"00000000000000000000111000000000" AFTER 08840 ns,
					"00000000000000000000000000000000" AFTER 08860 ns,
					"00000000000000000000111010000000" AFTER 08880 ns,
					"00000000000000000000000000000000" AFTER 08900 ns,
					"00000000000000000000111100000000" AFTER 08920 ns,
					"00000000000000000000000000000000" AFTER 08940 ns,
					"00000000000000000000111110000000" AFTER 08960 ns,
					"00000000000000000000000000000000" AFTER 08980 ns,
					"00000000000000000000000000000000" AFTER 09000 ns,
					"00000000000000000000000000000000" AFTER 09020 ns,
					"00000000000000000000000010000000" AFTER 09040 ns,
					"00000000000000000000000000000000" AFTER 09060 ns,
					"00000000000000000000000100000000" AFTER 09080 ns,
					"00000000000000000000000000000000" AFTER 09100 ns,
					"00000000000000000000000110000000" AFTER 09120 ns,
					"00000000000000000000000000000000" AFTER 09140 ns,
					"00000000000000000000001000000000" AFTER 09160 ns,
					"00000000000000000000000000000000" AFTER 09180 ns,
					"00000000000000000000001010000000" AFTER 09200 ns,
					"00000000000000000000000000000000" AFTER 09220 ns,
					"00000000000000000000001100000000" AFTER 09240 ns,
					"00000000000000000000000000000000" AFTER 09260 ns,
					"00000000000000000000001110000000" AFTER 09280 ns,
					"00000000000000000000000000000000" AFTER 09300 ns,
					"00000000000000000000010000000000" AFTER 09320 ns,
					"00000000000000000000000000000000" AFTER 09340 ns,
					"00000000000000000000010010000000" AFTER 09360 ns,
					"00000000000000000000000000000000" AFTER 09380 ns,
					"00000000000000000000010100000000" AFTER 09400 ns,
					"00000000000000000000000000000000" AFTER 09420 ns,
					"00000000000000000000010110000000" AFTER 09440 ns,
					"00000000000000000000000000000000" AFTER 09460 ns,
					"00000000000000000000011000000000" AFTER 09480 ns,
					"00000000000000000000000000000000" AFTER 09500 ns,
					"00000000000000000000011010000000" AFTER 09520 ns,
					"00000000000000000000000000000000" AFTER 09540 ns,
					"00000000000000000000011100000000" AFTER 09560 ns,
					"00000000000000000000000000000000" AFTER 09580 ns,
					"00000000000000000000011110000000" AFTER 09600 ns,
					"00000000000000000000000000000000" AFTER 09620 ns,
					"00000000000000000000100000000000" AFTER 09640 ns,
					"00000000000000000000000000000000" AFTER 09660 ns,
					"00000000000000000000100010000000" AFTER 09680 ns,
					"00000000000000000000000000000000" AFTER 09700 ns,
					"00000000000000000000100100000000" AFTER 09720 ns,
					"00000000000000000000000000000000" AFTER 09740 ns,
					"00000000000000000000100110000000" AFTER 09760 ns,
					"00000000000000000000000000000000" AFTER 09780 ns,
					"00000000000000000000101000000000" AFTER 09800 ns,
					"00000000000000000000000000000000" AFTER 09820 ns,
					"00000000000000000000101010000000" AFTER 09840 ns,
					"00000000000000000000000000000000" AFTER 09860 ns,
					"00000000000000000000101100000000" AFTER 09880 ns,
					"00000000000000000000000000000000" AFTER 09900 ns,
					"00000000000000000000101110000000" AFTER 09920 ns,
					"00000000000000000000000000000000" AFTER 09940 ns,
					"00000000000000000000110000000000" AFTER 09960 ns,
					"00000000000000000000000000000000" AFTER 09980 ns,
					"00000000000000000000110010000000" AFTER 10000 ns,
					"00000000000000000000000000000000" AFTER 10020 ns,
					"00000000000000000000110100000000" AFTER 10040 ns,
					"00000000000000000000000000000000" AFTER 10060 ns,
					"00000000000000000000110110000000" AFTER 10080 ns,
					"00000000000000000000000000000000" AFTER 10100 ns,
					"00000000000000000000111000000000" AFTER 10120 ns,
					"00000000000000000000000000000000" AFTER 10140 ns,
					"00000000000000000000111010000000" AFTER 10160 ns,
					"00000000000000000000000000000000" AFTER 10180 ns,
					"00000000000000000000111100000000" AFTER 10200 ns,
					"00000000000000000000000000000000" AFTER 10220 ns,
					"00000000000000000000111110000000" AFTER 10240 ns,
					"00000000000000000000000000000000" AFTER 10260 ns,
					"00000000000000000000000000000000" AFTER 10280 ns,
					"00000000000000000000000000000000" AFTER 10300 ns,
					"00000000000000000000000010000000" AFTER 10320 ns,
					"00000000000000000000000000000000" AFTER 10340 ns,
					"00000000000000000000000100000000" AFTER 10360 ns,
					"00000000000000000000000000000000" AFTER 10380 ns,
					"00000000000000000000000110000000" AFTER 10400 ns,
					"00000000000000000000000000000000" AFTER 10420 ns,
					"00000000000000000000001000000000" AFTER 10440 ns,
					"00000000000000000000000000000000" AFTER 10460 ns,
					"00000000000000000000001010000000" AFTER 10480 ns,
					"00000000000000000000000000000000" AFTER 10500 ns,
					"00000000000000000000001100000000" AFTER 10520 ns,
					"00000000000000000000000000000000" AFTER 10540 ns,
					"00000000000000000000001110000000" AFTER 10560 ns,
					"00000000000000000000000000000000" AFTER 10580 ns,
					"00000000000000000000010000000000" AFTER 10600 ns,
					"00000000000000000000000000000000" AFTER 10620 ns,
					"00000000000000000000010010000000" AFTER 10640 ns,
					"00000000000000000000000000000000" AFTER 10660 ns,
					"00000000000000000000010100000000" AFTER 10680 ns,
					"00000000000000000000000000000000" AFTER 10700 ns,
					"00000000000000000000010110000000" AFTER 10720 ns,
					"00000000000000000000000000000000" AFTER 10740 ns,
					"00000000000000000000011000000000" AFTER 10760 ns,
					"00000000000000000000000000000000" AFTER 10780 ns,
					"00000000000000000000011010000000" AFTER 10800 ns,
					"00000000000000000000000000000000" AFTER 10820 ns,
					"00000000000000000000011100000000" AFTER 10840 ns,
					"00000000000000000000000000000000" AFTER 10860 ns,
					"00000000000000000000011110000000" AFTER 10880 ns,
					"00000000000000000000000000000000" AFTER 10900 ns,
					"00000000000000000000100000000000" AFTER 10920 ns,
					"00000000000000000000000000000000" AFTER 10940 ns,
					"00000000000000000000100010000000" AFTER 10960 ns,
					"00000000000000000000000000000000" AFTER 10980 ns,
					"00000000000000000000100100000000" AFTER 11000 ns,
					"00000000000000000000000000000000" AFTER 11020 ns,
					"00000000000000000000100110000000" AFTER 11040 ns,
					"00000000000000000000000000000000" AFTER 11060 ns,
					"00000000000000000000101000000000" AFTER 11080 ns,
					"00000000000000000000000000000000" AFTER 11100 ns,
					"00000000000000000000101010000000" AFTER 11120 ns,
					"00000000000000000000000000000000" AFTER 11140 ns,
					"00000000000000000000101100000000" AFTER 11160 ns,
					"00000000000000000000000000000000" AFTER 11180 ns,
					"00000000000000000000101110000000" AFTER 11200 ns,
					"00000000000000000000000000000000" AFTER 11220 ns,
					"00000000000000000000110000000000" AFTER 11240 ns,
					"00000000000000000000000000000000" AFTER 11260 ns,
					"00000000000000000000110010000000" AFTER 11280 ns,
					"00000000000000000000000000000000" AFTER 11300 ns,
					"00000000000000000000110100000000" AFTER 11320 ns,
					"00000000000000000000000000000000" AFTER 11340 ns,
					"00000000000000000000110110000000" AFTER 11360 ns,
					"00000000000000000000000000000000" AFTER 11380 ns,
					"00000000000000000000111000000000" AFTER 11400 ns,
					"00000000000000000000000000000000" AFTER 11420 ns,
					"00000000000000000000111010000000" AFTER 11440 ns,
					"00000000000000000000000000000000" AFTER 11460 ns,
					"00000000000000000000111100000000" AFTER 11480 ns,
					"00000000000000000000000000000000" AFTER 11500 ns,
					"00000000000000000000111110000000" AFTER 11520 ns,
					"00000000000000000000000000000000" AFTER 11540 ns,
					"00000000000000000000000000000000" AFTER 11560 ns,
					"00000000000000000000000000000000" AFTER 11580 ns,
					"00000000000000000000000010000000" AFTER 11600 ns,
					"00000000000000000000000000000000" AFTER 11620 ns,
					"00000000000000000000000100000000" AFTER 11640 ns,
					"00000000000000000000000000000000" AFTER 11660 ns,
					"00000000000000000000000110000000" AFTER 11680 ns,
					"00000000000000000000000000000000" AFTER 11700 ns,
					"00000000000000000000001000000000" AFTER 11720 ns,
					"00000000000000000000000000000000" AFTER 11740 ns,
					"00000000000000000000001010000000" AFTER 11760 ns,
					"00000000000000000000000000000000" AFTER 11780 ns,
					"00000000000000000000001100000000" AFTER 11800 ns,
					"00000000000000000000000000000000" AFTER 11820 ns,
					"00000000000000000000001110000000" AFTER 11840 ns,
					"00000000000000000000000000000000" AFTER 11860 ns,
					"00000000000000000000010000000000" AFTER 11880 ns,
					"00000000000000000000000000000000" AFTER 11900 ns,
					"00000000000000000000010010000000" AFTER 11920 ns,
					"00000000000000000000000000000000" AFTER 11940 ns,
					"00000000000000000000010100000000" AFTER 11960 ns,
					"00000000000000000000000000000000" AFTER 11980 ns,
					"00000000000000000000010110000000" AFTER 12000 ns,
					"00000000000000000000000000000000" AFTER 12020 ns,
					"00000000000000000000011000000000" AFTER 12040 ns,
					"00000000000000000000000000000000" AFTER 12060 ns,
					"00000000000000000000011010000000" AFTER 12080 ns,
					"00000000000000000000000000000000" AFTER 12100 ns,
					"00000000000000000000011100000000" AFTER 12120 ns,
					"00000000000000000000000000000000" AFTER 12140 ns,
					"00000000000000000000011110000000" AFTER 12160 ns,
					"00000000000000000000000000000000" AFTER 12180 ns,
					"00000000000000000000100000000000" AFTER 12200 ns,
					"00000000000000000000000000000000" AFTER 12220 ns,
					"00000000000000000000100010000000" AFTER 12240 ns,
					"00000000000000000000000000000000" AFTER 12260 ns,
					"00000000000000000000100100000000" AFTER 12280 ns,
					"00000000000000000000000000000000" AFTER 12300 ns,
					"00000000000000000000100110000000" AFTER 12320 ns,
					"00000000000000000000000000000000" AFTER 12340 ns,
					"00000000000000000000101000000000" AFTER 12360 ns,
					"00000000000000000000000000000000" AFTER 12380 ns,
					"00000000000000000000101010000000" AFTER 12400 ns,
					"00000000000000000000000000000000" AFTER 12420 ns,
					"00000000000000000000101100000000" AFTER 12440 ns,
					"00000000000000000000000000000000" AFTER 12460 ns,
					"00000000000000000000101110000000" AFTER 12480 ns,
					"00000000000000000000000000000000" AFTER 12500 ns,
					"00000000000000000000110000000000" AFTER 12520 ns,
					"00000000000000000000000000000000" AFTER 12540 ns,
					"00000000000000000000110010000000" AFTER 12560 ns,
					"00000000000000000000000000000000" AFTER 12580 ns,
					"00000000000000000000110100000000" AFTER 12600 ns,
					"00000000000000000000000000000000" AFTER 12620 ns,
					"00000000000000000000110110000000" AFTER 12640 ns,
					"00000000000000000000000000000000" AFTER 12660 ns,
					"00000000000000000000111000000000" AFTER 12680 ns,
					"00000000000000000000000000000000" AFTER 12700 ns,
					"00000000000000000000111010000000" AFTER 12720 ns,
					"00000000000000000000000000000000" AFTER 12740 ns,
					"00000000000000000000111100000000" AFTER 12760 ns,
					"00000000000000000000000000000000" AFTER 12780 ns,
					"00000000000000000000111110000000" AFTER 12800 ns,
					"00000000000000000000000000000000" AFTER 12820 ns,
					"00000000000000000000000000000000" AFTER 12840 ns,
					"00000000000000000000000000000000" AFTER 12860 ns,
					"00000000000100000000000000000000" AFTER 12880 ns,
					"00000000000000000000000000000000" AFTER 12900 ns,
					"00000000001000000000000000000000" AFTER 12920 ns,
					"00000000000000000000000000000000" AFTER 12940 ns,
					"00000000001100000000000000000000" AFTER 12960 ns,
					"00000000000000000000000000000000" AFTER 12980 ns,
					"00000000010000000000000000000000" AFTER 13000 ns,
					"00000000000000000000000000000000" AFTER 13020 ns,
					"00000000010100000000000000000000" AFTER 13040 ns,
					"00000000000000000000000000000000" AFTER 13060 ns,
					"00000000011000000000000000000000" AFTER 13080 ns,
					"00000000000000000000000000000000" AFTER 13100 ns,
					"00000000011100000000000000000000" AFTER 13120 ns,
					"00000000000000000000000000000000" AFTER 13140 ns,
					"00000000100000000000000000000000" AFTER 13160 ns,
					"00000000000000000000000000000000" AFTER 13180 ns,
					"00000000100100000000000000000000" AFTER 13200 ns,
					"00000000000000000000000000000000" AFTER 13220 ns,
					"00000000101000000000000000000000" AFTER 13240 ns,
					"00000000000000000000000000000000" AFTER 13260 ns,
					"00000000101100000000000000000000" AFTER 13280 ns,
					"00000000000000000000000000000000" AFTER 13300 ns,
					"00000000110000000000000000000000" AFTER 13320 ns,
					"00000000000000000000000000000000" AFTER 13340 ns,
					"00000000110100000000000000000000" AFTER 13360 ns,
					"00000000000000000000000000000000" AFTER 13380 ns,
					"00000000111000000000000000000000" AFTER 13400 ns,
					"00000000000000000000000000000000" AFTER 13420 ns,
					"00000000111100000000000000000000" AFTER 13440 ns,
					"00000000000000000000000000000000" AFTER 13460 ns,
					"00000001000000000000000000000000" AFTER 13480 ns,
					"00000000000000000000000000000000" AFTER 13500 ns,
					"00000001000100000000000000000000" AFTER 13520 ns,
					"00000000000000000000000000000000" AFTER 13540 ns,
					"00000001001000000000000000000000" AFTER 13560 ns,
					"00000000000000000000000000000000" AFTER 13580 ns,
					"00000001001100000000000000000000" AFTER 13600 ns,
					"00000000000000000000000000000000" AFTER 13620 ns,
					"00000001010000000000000000000000" AFTER 13640 ns,
					"00000000000000000000000000000000" AFTER 13660 ns,
					"00000001010100000000000000000000" AFTER 13680 ns,
					"00000000000000000000000000000000" AFTER 13700 ns,
					"00000001011000000000000000000000" AFTER 13720 ns,
					"00000000000000000000000000000000" AFTER 13740 ns,
					"00000001011100000000000000000000" AFTER 13760 ns,
					"00000000000000000000000000000000" AFTER 13780 ns,
					"00000001100000000000000000000000" AFTER 13800 ns,
					"00000000000000000000000000000000" AFTER 13820 ns,
					"00000001100100000000000000000000" AFTER 13840 ns,
					"00000000000000000000000000000000" AFTER 13860 ns,
					"00000001101000000000000000000000" AFTER 13880 ns,
					"00000000000000000000000000000000" AFTER 13900 ns,
					"00000001101100000000000000000000" AFTER 13920 ns,
					"00000000000000000000000000000000" AFTER 13940 ns,
					"00000001110000000000000000000000" AFTER 13960 ns,
					"00000000000000000000000000000000" AFTER 13980 ns,
					"00000001110100000000000000000000" AFTER 14000 ns,
					"00000000000000000000000000000000" AFTER 14020 ns,
					"00000001111000000000000000000000" AFTER 14040 ns,
					"00000000000000000000000000000000" AFTER 14060 ns,
					"00000001111100000000000000000000" AFTER 14080 ns,
					"00000000000000000000000000000000" AFTER 14100 ns,
					"00000000000000000000000000000000" AFTER 14120 ns,
					"00000000000000000000000000000000" AFTER 14140 ns,
					"00000000000100000000000000000000" AFTER 14160 ns,
					"00000000000000000000000000000000" AFTER 14180 ns,
					"00000000001000000000000000000000" AFTER 14200 ns,
					"00000000000000000000000000000000" AFTER 14220 ns,
					"00000000001100000000000000000000" AFTER 14240 ns,
					"00000000000000000000000000000000" AFTER 14260 ns,
					"00000000010000000000000000000000" AFTER 14280 ns,
					"00000000000000000000000000000000" AFTER 14300 ns,
					"00000000010100000000000000000000" AFTER 14320 ns,
					"00000000000000000000000000000000" AFTER 14340 ns,
					"00000000011000000000000000000000" AFTER 14360 ns,
					"00000000000000000000000000000000" AFTER 14380 ns,
					"00000000011100000000000000000000" AFTER 14400 ns,
					"00000000000000000000000000000000" AFTER 14420 ns,
					"00000000100000000000000000000000" AFTER 14440 ns,
					"00000000000000000000000000000000" AFTER 14460 ns,
					"00000000100100000000000000000000" AFTER 14480 ns,
					"00000000000000000000000000000000" AFTER 14500 ns,
					"00000000101000000000000000000000" AFTER 14520 ns,
					"00000000000000000000000000000000" AFTER 14540 ns,
					"00000000101100000000000000000000" AFTER 14560 ns,
					"00000000000000000000000000000000" AFTER 14580 ns,
					"00000000110000000000000000000000" AFTER 14600 ns,
					"00000000000000000000000000000000" AFTER 14620 ns,
					"00000000110100000000000000000000" AFTER 14640 ns,
					"00000000000000000000000000000000" AFTER 14660 ns,
					"00000000111000000000000000000000" AFTER 14680 ns,
					"00000000000000000000000000000000" AFTER 14700 ns,
					"00000000111100000000000000000000" AFTER 14720 ns,
					"00000000000000000000000000000000" AFTER 14740 ns,
					"00000001000000000000000000000000" AFTER 14760 ns,
					"00000000000000000000000000000000" AFTER 14780 ns,
					"00000001000100000000000000000000" AFTER 14800 ns,
					"00000000000000000000000000000000" AFTER 14820 ns,
					"00000001001000000000000000000000" AFTER 14840 ns,
					"00000000000000000000000000000000" AFTER 14860 ns,
					"00000001001100000000000000000000" AFTER 14880 ns,
					"00000000000000000000000000000000" AFTER 14900 ns,
					"00000001010000000000000000000000" AFTER 14920 ns,
					"00000000000000000000000000000000" AFTER 14940 ns,
					"00000001010100000000000000000000" AFTER 14960 ns,
					"00000000000000000000000000000000" AFTER 14980 ns,
					"00000001011000000000000000000000" AFTER 15000 ns,
					"00000000000000000000000000000000" AFTER 15020 ns,
					"00000001011100000000000000000000" AFTER 15040 ns,
					"00000000000000000000000000000000" AFTER 15060 ns,
					"00000001100000000000000000000000" AFTER 15080 ns,
					"00000000000000000000000000000000" AFTER 15100 ns,
					"00000001100100000000000000000000" AFTER 15120 ns,
					"00000000000000000000000000000000" AFTER 15140 ns,
					"00000001101000000000000000000000" AFTER 15160 ns,
					"00000000000000000000000000000000" AFTER 15180 ns,
					"00000001101100000000000000000000" AFTER 15200 ns,
					"00000000000000000000000000000000" AFTER 15220 ns,
					"00000001110000000000000000000000" AFTER 15240 ns,
					"00000000000000000000000000000000" AFTER 15260 ns,
					"00000001110100000000000000000000" AFTER 15280 ns,
					"00000000000000000000000000000000" AFTER 15300 ns,
					"00000001111000000000000000000000" AFTER 15320 ns,
					"00000000000000000000000000000000" AFTER 15340 ns,
					"00000001111100000000000000000000" AFTER 15360 ns,
					"00000000000000000000000000000000" AFTER 15380 ns,
					"00000000000000000000000000000000" AFTER 15400 ns,
					"00000000000000000000000000000000" AFTER 15420 ns,
					"00000000000100000000000000000000" AFTER 15440 ns,
					"00000000000000000000000000000000" AFTER 15460 ns,
					"00000000001000000000000000000000" AFTER 15480 ns,
					"00000000000000000000000000000000" AFTER 15500 ns,
					"00000000001100000000000000000000" AFTER 15520 ns,
					"00000000000000000000000000000000" AFTER 15540 ns,
					"00000000010000000000000000000000" AFTER 15560 ns,
					"00000000000000000000000000000000" AFTER 15580 ns,
					"00000000010100000000000000000000" AFTER 15600 ns,
					"00000000000000000000000000000000" AFTER 15620 ns,
					"00000000011000000000000000000000" AFTER 15640 ns,
					"00000000000000000000000000000000" AFTER 15660 ns,
					"00000000011100000000000000000000" AFTER 15680 ns,
					"00000000000000000000000000000000" AFTER 15700 ns,
					"00000000100000000000000000000000" AFTER 15720 ns,
					"00000000000000000000000000000000" AFTER 15740 ns,
					"00000000100100000000000000000000" AFTER 15760 ns,
					"00000000000000000000000000000000" AFTER 15780 ns,
					"00000000101000000000000000000000" AFTER 15800 ns,
					"00000000000000000000000000000000" AFTER 15820 ns,
					"00000000101100000000000000000000" AFTER 15840 ns,
					"00000000000000000000000000000000" AFTER 15860 ns,
					"00000000110000000000000000000000" AFTER 15880 ns,
					"00000000000000000000000000000000" AFTER 15900 ns,
					"00000000110100000000000000000000" AFTER 15920 ns,
					"00000000000000000000000000000000" AFTER 15940 ns,
					"00000000111000000000000000000000" AFTER 15960 ns,
					"00000000000000000000000000000000" AFTER 15980 ns,
					"00000000111100000000000000000000" AFTER 16000 ns,
					"00000000000000000000000000000000" AFTER 16020 ns,
					"00000001000000000000000000000000" AFTER 16040 ns,
					"00000000000000000000000000000000" AFTER 16060 ns,
					"00000001000100000000000000000000" AFTER 16080 ns,
					"00000000000000000000000000000000" AFTER 16100 ns,
					"00000001001000000000000000000000" AFTER 16120 ns,
					"00000000000000000000000000000000" AFTER 16140 ns,
					"00000001001100000000000000000000" AFTER 16160 ns,
					"00000000000000000000000000000000" AFTER 16180 ns,
					"00000001010000000000000000000000" AFTER 16200 ns,
					"00000000000000000000000000000000" AFTER 16220 ns,
					"00000001010100000000000000000000" AFTER 16240 ns,
					"00000000000000000000000000000000" AFTER 16260 ns,
					"00000001011000000000000000000000" AFTER 16280 ns,
					"00000000000000000000000000000000" AFTER 16300 ns,
					"00000001011100000000000000000000" AFTER 16320 ns,
					"00000000000000000000000000000000" AFTER 16340 ns,
					"00000001100000000000000000000000" AFTER 16360 ns,
					"00000000000000000000000000000000" AFTER 16380 ns,
					"00000001100100000000000000000000" AFTER 16400 ns,
					"00000000000000000000000000000000" AFTER 16420 ns,
					"00000001101000000000000000000000" AFTER 16440 ns,
					"00000000000000000000000000000000" AFTER 16460 ns,
					"00000001101100000000000000000000" AFTER 16480 ns,
					"00000000000000000000000000000000" AFTER 16500 ns,
					"00000001110000000000000000000000" AFTER 16520 ns,
					"00000000000000000000000000000000" AFTER 16540 ns,
					"00000001110100000000000000000000" AFTER 16560 ns,
					"00000000000000000000000000000000" AFTER 16580 ns,
					"00000001111000000000000000000000" AFTER 16600 ns,
					"00000000000000000000000000000000" AFTER 16620 ns,
					"00000001111100000000000000000000" AFTER 16640 ns,
					"00000000000000000000000000000000" AFTER 16660 ns,
					"00000000000000000000000000000000" AFTER 16680 ns,
					"00000000000000000000000000000000" AFTER 16700 ns,
					"00000000000000000000000010000000" AFTER 16720 ns,
					"00000000000000000000000000000000" AFTER 16740 ns,
					"00000000000000000000000100000000" AFTER 16760 ns,
					"00000000000000000000000000000000" AFTER 16780 ns,
					"00000000000000000000000110000000" AFTER 16800 ns,
					"00000000000000000000000000000000" AFTER 16820 ns,
					"00000000000000000000001000000000" AFTER 16840 ns,
					"00000000000000000000000000000000" AFTER 16860 ns,
					"00000000000000000000001010000000" AFTER 16880 ns,
					"00000000000000000000000000000000" AFTER 16900 ns,
					"00000000000000000000001100000000" AFTER 16920 ns,
					"00000000000000000000000000000000" AFTER 16940 ns,
					"00000000000000000000001110000000" AFTER 16960 ns,
					"00000000000000000000000000000000" AFTER 16980 ns,
					"00000000000000000000010000000000" AFTER 17000 ns,
					"00000000000000000000000000000000" AFTER 17020 ns,
					"00000000000000000000010010000000" AFTER 17040 ns,
					"00000000000000000000000000000000" AFTER 17060 ns,
					"00000000000000000000010100000000" AFTER 17080 ns,
					"00000000000000000000000000000000" AFTER 17100 ns,
					"00000000000000000000010110000000" AFTER 17120 ns,
					"00000000000000000000000000000000" AFTER 17140 ns,
					"00000000000000000000011000000000" AFTER 17160 ns,
					"00000000000000000000000000000000" AFTER 17180 ns,
					"00000000000000000000011010000000" AFTER 17200 ns,
					"00000000000000000000000000000000" AFTER 17220 ns,
					"00000000000000000000011100000000" AFTER 17240 ns,
					"00000000000000000000000000000000" AFTER 17260 ns,
					"00000000000000000000011110000000" AFTER 17280 ns,
					"00000000000000000000000000000000" AFTER 17300 ns,
					"00000000000000000000100000000000" AFTER 17320 ns,
					"00000000000000000000000000000000" AFTER 17340 ns,
					"00000000000000000000100010000000" AFTER 17360 ns,
					"00000000000000000000000000000000" AFTER 17380 ns,
					"00000000000000000000100100000000" AFTER 17400 ns,
					"00000000000000000000000000000000" AFTER 17420 ns,
					"00000000000000000000100110000000" AFTER 17440 ns,
					"00000000000000000000000000000000" AFTER 17460 ns,
					"00000000000000000000101000000000" AFTER 17480 ns,
					"00000000000000000000000000000000" AFTER 17500 ns,
					"00000000000000000000101010000000" AFTER 17520 ns,
					"00000000000000000000000000000000" AFTER 17540 ns,
					"00000000000000000000101100000000" AFTER 17560 ns,
					"00000000000000000000000000000000" AFTER 17580 ns,
					"00000000000000000000101110000000" AFTER 17600 ns,
					"00000000000000000000000000000000" AFTER 17620 ns,
					"00000000000000000000110000000000" AFTER 17640 ns,
					"00000000000000000000000000000000" AFTER 17660 ns,
					"00000000000000000000110010000000" AFTER 17680 ns,
					"00000000000000000000000000000000" AFTER 17700 ns,
					"00000000000000000000110100000000" AFTER 17720 ns,
					"00000000000000000000000000000000" AFTER 17740 ns,
					"00000000000000000000110110000000" AFTER 17760 ns,
					"00000000000000000000000000000000" AFTER 17780 ns,
					"00000000000000000000111000000000" AFTER 17800 ns,
					"00000000000000000000000000000000" AFTER 17820 ns,
					"00000000000000000000111010000000" AFTER 17840 ns,
					"00000000000000000000000000000000" AFTER 17860 ns,
					"00000000000000000000111100000000" AFTER 17880 ns,
					"00000000000000000000000000000000" AFTER 17900 ns,
					"00000000000000000000111110000000" AFTER 17920 ns,
					"00000000000000000000000000000000" AFTER 17940 ns,
					"00000000000000000000000000000000" AFTER 17960 ns,
					"00000000000000000000000000000000" AFTER 17980 ns,
					"00000000000000000000000010000000" AFTER 18000 ns,
					"00000000000000000000000000000000" AFTER 18020 ns,
					"00000000000000000000000100000000" AFTER 18040 ns,
					"00000000000000000000000000000000" AFTER 18060 ns,
					"00000000000000000000000110000000" AFTER 18080 ns,
					"00000000000000000000000000000000" AFTER 18100 ns,
					"00000000000000000000001000000000" AFTER 18120 ns,
					"00000000000000000000000000000000" AFTER 18140 ns,
					"00000000000000000000001010000000" AFTER 18160 ns,
					"00000000000000000000000000000000" AFTER 18180 ns,
					"00000000000000000000001100000000" AFTER 18200 ns,
					"00000000000000000000000000000000" AFTER 18220 ns,
					"00000000000000000000001110000000" AFTER 18240 ns,
					"00000000000000000000000000000000" AFTER 18260 ns,
					"00000000000000000000010000000000" AFTER 18280 ns,
					"00000000000000000000000000000000" AFTER 18300 ns,
					"00000000000000000000010010000000" AFTER 18320 ns,
					"00000000000000000000000000000000" AFTER 18340 ns,
					"00000000000000000000010100000000" AFTER 18360 ns,
					"00000000000000000000000000000000" AFTER 18380 ns,
					"00000000000000000000010110000000" AFTER 18400 ns,
					"00000000000000000000000000000000" AFTER 18420 ns,
					"00000000000000000000011000000000" AFTER 18440 ns,
					"00000000000000000000000000000000" AFTER 18460 ns,
					"00000000000000000000011010000000" AFTER 18480 ns,
					"00000000000000000000000000000000" AFTER 18500 ns,
					"00000000000000000000011100000000" AFTER 18520 ns,
					"00000000000000000000000000000000" AFTER 18540 ns,
					"00000000000000000000011110000000" AFTER 18560 ns,
					"00000000000000000000000000000000" AFTER 18580 ns,
					"00000000000000000000100000000000" AFTER 18600 ns,
					"00000000000000000000000000000000" AFTER 18620 ns,
					"00000000000000000000100010000000" AFTER 18640 ns,
					"00000000000000000000000000000000" AFTER 18660 ns,
					"00000000000000000000100100000000" AFTER 18680 ns,
					"00000000000000000000000000000000" AFTER 18700 ns,
					"00000000000000000000100110000000" AFTER 18720 ns,
					"00000000000000000000000000000000" AFTER 18740 ns,
					"00000000000000000000101000000000" AFTER 18760 ns,
					"00000000000000000000000000000000" AFTER 18780 ns,
					"00000000000000000000101010000000" AFTER 18800 ns,
					"00000000000000000000000000000000" AFTER 18820 ns,
					"00000000000000000000101100000000" AFTER 18840 ns,
					"00000000000000000000000000000000" AFTER 18860 ns,
					"00000000000000000000101110000000" AFTER 18880 ns,
					"00000000000000000000000000000000" AFTER 18900 ns,
					"00000000000000000000110000000000" AFTER 18920 ns,
					"00000000000000000000000000000000" AFTER 18940 ns,
					"00000000000000000000110010000000" AFTER 18960 ns,
					"00000000000000000000000000000000" AFTER 18980 ns,
					"00000000000000000000110100000000" AFTER 19000 ns,
					"00000000000000000000000000000000" AFTER 19020 ns,
					"00000000000000000000110110000000" AFTER 19040 ns,
					"00000000000000000000000000000000" AFTER 19060 ns,
					"00000000000000000000111000000000" AFTER 19080 ns,
					"00000000000000000000000000000000" AFTER 19100 ns,
					"00000000000000000000111010000000" AFTER 19120 ns,
					"00000000000000000000000000000000" AFTER 19140 ns,
					"00000000000000000000111100000000" AFTER 19160 ns,
					"00000000000000000000000000000000" AFTER 19180 ns,
					"00000000000000000000111110000000" AFTER 19200 ns,
					"00000000000000000000000000000000" AFTER 19220 ns,
					"00000000000000000000000000000000" AFTER 19240 ns,
					"00000000000000000000000000000000" AFTER 19260 ns,
					"00000000000000000000000010000000" AFTER 19280 ns,
					"00000000000000000000000000000000" AFTER 19300 ns,
					"00000000000000000000000100000000" AFTER 19320 ns,
					"00000000000000000000000000000000" AFTER 19340 ns,
					"00000000000000000000000110000000" AFTER 19360 ns,
					"00000000000000000000000000000000" AFTER 19380 ns,
					"00000000000000000000001000000000" AFTER 19400 ns,
					"00000000000000000000000000000000" AFTER 19420 ns,
					"00000000000000000000001010000000" AFTER 19440 ns,
					"00000000000000000000000000000000" AFTER 19460 ns,
					"00000000000000000000001100000000" AFTER 19480 ns,
					"00000000000000000000000000000000" AFTER 19500 ns,
					"00000000000000000000001110000000" AFTER 19520 ns,
					"00000000000000000000000000000000" AFTER 19540 ns,
					"00000000000000000000010000000000" AFTER 19560 ns,
					"00000000000000000000000000000000" AFTER 19580 ns,
					"00000000000000000000010010000000" AFTER 19600 ns,
					"00000000000000000000000000000000" AFTER 19620 ns,
					"00000000000000000000010100000000" AFTER 19640 ns,
					"00000000000000000000000000000000" AFTER 19660 ns,
					"00000000000000000000010110000000" AFTER 19680 ns,
					"00000000000000000000000000000000" AFTER 19700 ns,
					"00000000000000000000011000000000" AFTER 19720 ns,
					"00000000000000000000000000000000" AFTER 19740 ns,
					"00000000000000000000011010000000" AFTER 19760 ns,
					"00000000000000000000000000000000" AFTER 19780 ns,
					"00000000000000000000011100000000" AFTER 19800 ns,
					"00000000000000000000000000000000" AFTER 19820 ns,
					"00000000000000000000011110000000" AFTER 19840 ns,
					"00000000000000000000000000000000" AFTER 19860 ns,
					"00000000000000000000100000000000" AFTER 19880 ns,
					"00000000000000000000000000000000" AFTER 19900 ns,
					"00000000000000000000100010000000" AFTER 19920 ns,
					"00000000000000000000000000000000" AFTER 19940 ns,
					"00000000000000000000100100000000" AFTER 19960 ns,
					"00000000000000000000000000000000" AFTER 19980 ns,
					"00000000000000000000100110000000" AFTER 20000 ns,
					"00000000000000000000000000000000" AFTER 20020 ns,
					"00000000000000000000101000000000" AFTER 20040 ns,
					"00000000000000000000000000000000" AFTER 20060 ns,
					"00000000000000000000101010000000" AFTER 20080 ns,
					"00000000000000000000000000000000" AFTER 20100 ns,
					"00000000000000000000101100000000" AFTER 20120 ns,
					"00000000000000000000000000000000" AFTER 20140 ns,
					"00000000000000000000101110000000" AFTER 20160 ns,
					"00000000000000000000000000000000" AFTER 20180 ns,
					"00000000000000000000110000000000" AFTER 20200 ns,
					"00000000000000000000000000000000" AFTER 20220 ns,
					"00000000000000000000110010000000" AFTER 20240 ns,
					"00000000000000000000000000000000" AFTER 20260 ns,
					"00000000000000000000110100000000" AFTER 20280 ns,
					"00000000000000000000000000000000" AFTER 20300 ns,
					"00000000000000000000110110000000" AFTER 20320 ns,
					"00000000000000000000000000000000" AFTER 20340 ns,
					"00000000000000000000111000000000" AFTER 20360 ns,
					"00000000000000000000000000000000" AFTER 20380 ns,
					"00000000000000000000111010000000" AFTER 20400 ns,
					"00000000000000000000000000000000" AFTER 20420 ns,
					"00000000000000000000111100000000" AFTER 20440 ns,
					"00000000000000000000000000000000" AFTER 20460 ns,
					"00000000000000000000111110000000" AFTER 20480 ns,
					"00000000000000000000000000000000" AFTER 20500 ns,
					"00000000000000000000000000000000" AFTER 20520 ns,
					"00000000000000000000000000000000" AFTER 20540 ns,
					"00000000000000000000000010000000" AFTER 20560 ns,
					"00000000000000000000000000000000" AFTER 20580 ns,
					"00000000000000000000000100000000" AFTER 20600 ns,
					"00000000000000000000000000000000" AFTER 20620 ns,
					"00000000000000000000000110000000" AFTER 20640 ns,
					"00000000000000000000000000000000" AFTER 20660 ns,
					"00000000000000000000001000000000" AFTER 20680 ns,
					"00000000000000000000000000000000" AFTER 20700 ns,
					"00000000000000000000001010000000" AFTER 20720 ns,
					"00000000000000000000000000000000" AFTER 20740 ns,
					"00000000000000000000001100000000" AFTER 20760 ns,
					"00000000000000000000000000000000" AFTER 20780 ns,
					"00000000000000000000001110000000" AFTER 20800 ns,
					"00000000000000000000000000000000" AFTER 20820 ns,
					"00000000000000000000010000000000" AFTER 20840 ns,
					"00000000000000000000000000000000" AFTER 20860 ns,
					"00000000000000000000010010000000" AFTER 20880 ns,
					"00000000000000000000000000000000" AFTER 20900 ns,
					"00000000000000000000010100000000" AFTER 20920 ns,
					"00000000000000000000000000000000" AFTER 20940 ns,
					"00000000000000000000010110000000" AFTER 20960 ns,
					"00000000000000000000000000000000" AFTER 20980 ns,
					"00000000000000000000011000000000" AFTER 21000 ns,
					"00000000000000000000000000000000" AFTER 21020 ns,
					"00000000000000000000011010000000" AFTER 21040 ns,
					"00000000000000000000000000000000" AFTER 21060 ns,
					"00000000000000000000011100000000" AFTER 21080 ns,
					"00000000000000000000000000000000" AFTER 21100 ns,
					"00000000000000000000011110000000" AFTER 21120 ns,
					"00000000000000000000000000000000" AFTER 21140 ns,
					"00000000000000000000100000000000" AFTER 21160 ns,
					"00000000000000000000000000000000" AFTER 21180 ns,
					"00000000000000000000100010000000" AFTER 21200 ns,
					"00000000000000000000000000000000" AFTER 21220 ns,
					"00000000000000000000100100000000" AFTER 21240 ns,
					"00000000000000000000000000000000" AFTER 21260 ns,
					"00000000000000000000100110000000" AFTER 21280 ns,
					"00000000000000000000000000000000" AFTER 21300 ns,
					"00000000000000000000101000000000" AFTER 21320 ns,
					"00000000000000000000000000000000" AFTER 21340 ns,
					"00000000000000000000101010000000" AFTER 21360 ns,
					"00000000000000000000000000000000" AFTER 21380 ns,
					"00000000000000000000101100000000" AFTER 21400 ns,
					"00000000000000000000000000000000" AFTER 21420 ns,
					"00000000000000000000101110000000" AFTER 21440 ns,
					"00000000000000000000000000000000" AFTER 21460 ns,
					"00000000000000000000110000000000" AFTER 21480 ns,
					"00000000000000000000000000000000" AFTER 21500 ns,
					"00000000000000000000110010000000" AFTER 21520 ns,
					"00000000000000000000000000000000" AFTER 21540 ns,
					"00000000000000000000110100000000" AFTER 21560 ns,
					"00000000000000000000000000000000" AFTER 21580 ns,
					"00000000000000000000110110000000" AFTER 21600 ns,
					"00000000000000000000000000000000" AFTER 21620 ns,
					"00000000000000000000111000000000" AFTER 21640 ns,
					"00000000000000000000000000000000" AFTER 21660 ns,
					"00000000000000000000111010000000" AFTER 21680 ns,
					"00000000000000000000000000000000" AFTER 21700 ns,
					"00000000000000000000111100000000" AFTER 21720 ns,
					"00000000000000000000000000000000" AFTER 21740 ns,
					"00000000000000000000111110000000" AFTER 21760 ns,
					"00000000000000000000000000000000" AFTER 21780 ns,
					"00000000000011111000000000000000" AFTER 21800 ns,
					"00000000000000000000000000000000" AFTER 21820 ns,
					"00000000000011110000000010000000" AFTER 21840 ns,
					"00000000000000000000000000000000" AFTER 21860 ns,
					"00000000000011101000000100000000" AFTER 21880 ns,
					"00000000000000000000000000000000" AFTER 21900 ns,
					"00000000000011100000000110000000" AFTER 21920 ns,
					"00000000000000000000000000000000" AFTER 21940 ns,
					"00000000000011011000001000000000" AFTER 21960 ns,
					"00000000000000000000000000000000" AFTER 21980 ns,
					"00000000000011010000001010000000" AFTER 22000 ns,
					"00000000000000000000000000000000" AFTER 22020 ns,
					"00000000000011001000001100000000" AFTER 22040 ns,
					"00000000000000000000000000000000" AFTER 22060 ns,
					"00000000000011000000001110000000" AFTER 22080 ns,
					"00000000000000000000000000000000" AFTER 22100 ns,
					"00000000000010111000010000000000" AFTER 22120 ns,
					"00000000000000000000000000000000" AFTER 22140 ns,
					"00000000000010110000010010000000" AFTER 22160 ns,
					"00000000000000000000000000000000" AFTER 22180 ns,
					"00000000000010101000010100000000" AFTER 22200 ns,
					"00000000000000000000000000000000" AFTER 22220 ns,
					"00000000000010100000010110000000" AFTER 22240 ns,
					"00000000000000000000000000000000" AFTER 22260 ns,
					"00000000000010011000011000000000" AFTER 22280 ns,
					"00000000000000000000000000000000" AFTER 22300 ns,
					"00000000000010010000011010000000" AFTER 22320 ns,
					"00000000000000000000000000000000" AFTER 22340 ns,
					"00000000000010001000011100000000" AFTER 22360 ns,
					"00000000000000000000000000000000" AFTER 22380 ns,
					"00000000000010000000011110000000" AFTER 22400 ns,
					"00000000000000000000000000000000" AFTER 22420 ns,
					"00000000000001111000100000000000" AFTER 22440 ns,
					"00000000000000000000000000000000" AFTER 22460 ns,
					"00000000000001110000100010000000" AFTER 22480 ns,
					"00000000000000000000000000000000" AFTER 22500 ns,
					"00000000000001101000100100000000" AFTER 22520 ns,
					"00000000000000000000000000000000" AFTER 22540 ns,
					"00000000000001100000100110000000" AFTER 22560 ns,
					"00000000000000000000000000000000" AFTER 22580 ns,
					"00000000000001011000101000000000" AFTER 22600 ns,
					"00000000000000000000000000000000" AFTER 22620 ns,
					"00000000000001010000101010000000" AFTER 22640 ns,
					"00000000000000000000000000000000" AFTER 22660 ns,
					"00000000000001001000101100000000" AFTER 22680 ns,
					"00000000000000000000000000000000" AFTER 22700 ns,
					"00000000000001000000101110000000" AFTER 22720 ns,
					"00000000000000000000000000000000" AFTER 22740 ns,
					"00000000000000111000110000000000" AFTER 22760 ns,
					"00000000000000000000000000000000" AFTER 22780 ns,
					"00000000000000110000110010000000" AFTER 22800 ns,
					"00000000000000000000000000000000" AFTER 22820 ns,
					"00000000000000101000110100000000" AFTER 22840 ns,
					"00000000000000000000000000000000" AFTER 22860 ns,
					"00000000000000100000110110000000" AFTER 22880 ns,
					"00000000000000000000000000000000" AFTER 22900 ns,
					"00000000000000011000111000000000" AFTER 22920 ns,
					"00000000000000000000000000000000" AFTER 22940 ns,
					"00000000000000010000111010000000" AFTER 22960 ns,
					"00000000000000000000000000000000" AFTER 22980 ns,
					"00000000000000001000111100000000" AFTER 23000 ns,
					"00000000000000000000000000000000" AFTER 23020 ns,
					"00000000000000000000111110000000" AFTER 23040 ns,
					"00000000000000000000000000000000" AFTER 23060 ns,
					"00000000000011111000000000000000" AFTER 23080 ns,
					"00000000000000000000000000000000" AFTER 23100 ns,
					"00000000000111110000000010000000" AFTER 23120 ns,
					"00000000000000000000000000000000" AFTER 23140 ns,
					"00000000001011101000000100000000" AFTER 23160 ns,
					"00000000000000000000000000000000" AFTER 23180 ns,
					"00000000001111100000000110000000" AFTER 23200 ns,
					"00000000000000000000000000000000" AFTER 23220 ns,
					"00000000010011011000001000000000" AFTER 23240 ns,
					"00000000000000000000000000000000" AFTER 23260 ns,
					"00000000010111010000001010000000" AFTER 23280 ns,
					"00000000000000000000000000000000" AFTER 23300 ns,
					"00000000011011001000001100000000" AFTER 23320 ns,
					"00000000000000000000000000000000" AFTER 23340 ns,
					"00000000011111000000001110000000" AFTER 23360 ns,
					"00000000000000000000000000000000" AFTER 23380 ns,
					"00000000100010111000010000000000" AFTER 23400 ns,
					"00000000000000000000000000000000" AFTER 23420 ns,
					"00000000100110110000010010000000" AFTER 23440 ns,
					"00000000000000000000000000000000" AFTER 23460 ns,
					"00000000101010101000010100000000" AFTER 23480 ns,
					"00000000000000000000000000000000" AFTER 23500 ns,
					"00000000101110100000010110000000" AFTER 23520 ns,
					"00000000000000000000000000000000" AFTER 23540 ns,
					"00000000110010011000011000000000" AFTER 23560 ns,
					"00000000000000000000000000000000" AFTER 23580 ns,
					"00000000110110010000011010000000" AFTER 23600 ns,
					"00000000000000000000000000000000" AFTER 23620 ns,
					"00000000111010001000011100000000" AFTER 23640 ns,
					"00000000000000000000000000000000" AFTER 23660 ns,
					"00000000111110000000011110000000" AFTER 23680 ns,
					"00000000000000000000000000000000" AFTER 23700 ns,
					"00000001000001111000100000000000" AFTER 23720 ns,
					"00000000000000000000000000000000" AFTER 23740 ns,
					"00000001000101110000100010000000" AFTER 23760 ns,
					"00000000000000000000000000000000" AFTER 23780 ns,
					"00000001001001101000100100000000" AFTER 23800 ns,
					"00000000000000000000000000000000" AFTER 23820 ns,
					"00000001001101100000100110000000" AFTER 23840 ns,
					"00000000000000000000000000000000" AFTER 23860 ns,
					"00000001010001011000101000000000" AFTER 23880 ns,
					"00000000000000000000000000000000" AFTER 23900 ns,
					"00000001010101010000101010000000" AFTER 23920 ns,
					"00000000000000000000000000000000" AFTER 23940 ns,
					"00000001011001001000101100000000" AFTER 23960 ns,
					"00000000000000000000000000000000" AFTER 23980 ns,
					"00000001011101000000101110000000" AFTER 24000 ns,
					"00000000000000000000000000000000" AFTER 24020 ns,
					"00000001100000111000110000000000" AFTER 24040 ns,
					"00000000000000000000000000000000" AFTER 24060 ns,
					"00000001100100110000110010000000" AFTER 24080 ns,
					"00000000000000000000000000000000" AFTER 24100 ns,
					"00000001101000101000110100000000" AFTER 24120 ns,
					"00000000000000000000000000000000" AFTER 24140 ns,
					"00000001101100100000110110000000" AFTER 24160 ns,
					"00000000000000000000000000000000" AFTER 24180 ns,
					"00000001110000011000111000000000" AFTER 24200 ns,
					"00000000000000000000000000000000" AFTER 24220 ns,
					"00000001110100010000111010000000" AFTER 24240 ns,
					"00000000000000000000000000000000" AFTER 24260 ns,
					"00000001111000001000111100000000" AFTER 24280 ns,
					"00000000000000000000000000000000" AFTER 24300 ns,
					"00000001111100000000111110000000" AFTER 24320 ns,
					"00000000000000000000000000000000" AFTER 24340 ns,
					"00000000000000000000000000000000" AFTER 24360 ns,
					"00000000000000000000000000000000" AFTER 24380 ns,
					"00000000000000000000000010000000" AFTER 24400 ns,
					"00000000000000000000000000000000" AFTER 24420 ns,
					"00000000000000000000000100000000" AFTER 24440 ns,
					"00000000000000000000000000000000" AFTER 24460 ns,
					"00000000000000000000000110000000" AFTER 24480 ns,
					"00000000000000000000000000000000" AFTER 24500 ns,
					"00000000000000000000001000000000" AFTER 24520 ns,
					"00000000000000000000000000000000" AFTER 24540 ns,
					"00000000000000000000001010000000" AFTER 24560 ns,
					"00000000000000000000000000000000" AFTER 24580 ns,
					"00000000000000000000001100000000" AFTER 24600 ns,
					"00000000000000000000000000000000" AFTER 24620 ns,
					"00000000000000000000001110000000" AFTER 24640 ns,
					"00000000000000000000000000000000" AFTER 24660 ns,
					"00000000000000000000010000000000" AFTER 24680 ns,
					"00000000000000000000000000000000" AFTER 24700 ns,
					"00000000000000000000010010000000" AFTER 24720 ns,
					"00000000000000000000000000000000" AFTER 24740 ns,
					"00000000000000000000010100000000" AFTER 24760 ns,
					"00000000000000000000000000000000" AFTER 24780 ns,
					"00000000000000000000010110000000" AFTER 24800 ns,
					"00000000000000000000000000000000" AFTER 24820 ns,
					"00000000000000000000011000000000" AFTER 24840 ns,
					"00000000000000000000000000000000" AFTER 24860 ns,
					"00000000000000000000011010000000" AFTER 24880 ns,
					"00000000000000000000000000000000" AFTER 24900 ns,
					"00000000000000000000011100000000" AFTER 24920 ns,
					"00000000000000000000000000000000" AFTER 24940 ns,
					"00000000000000000000011110000000" AFTER 24960 ns,
					"00000000000000000000000000000000" AFTER 24980 ns,
					"00000000000000000000100000000000" AFTER 25000 ns,
					"00000000000000000000000000000000" AFTER 25020 ns,
					"00000000000000000000100010000000" AFTER 25040 ns,
					"00000000000000000000000000000000" AFTER 25060 ns,
					"00000000000000000000100100000000" AFTER 25080 ns,
					"00000000000000000000000000000000" AFTER 25100 ns,
					"00000000000000000000100110000000" AFTER 25120 ns,
					"00000000000000000000000000000000" AFTER 25140 ns,
					"00000000000000000000101000000000" AFTER 25160 ns,
					"00000000000000000000000000000000" AFTER 25180 ns,
					"00000000000000000000101010000000" AFTER 25200 ns,
					"00000000000000000000000000000000" AFTER 25220 ns,
					"00000000000000000000101100000000" AFTER 25240 ns,
					"00000000000000000000000000000000" AFTER 25260 ns,
					"00000000000000000000101110000000" AFTER 25280 ns,
					"00000000000000000000000000000000" AFTER 25300 ns,
					"00000000000000000000110000000000" AFTER 25320 ns,
					"00000000000000000000000000000000" AFTER 25340 ns,
					"00000000000000000000110010000000" AFTER 25360 ns,
					"00000000000000000000000000000000" AFTER 25380 ns,
					"00000000000000000000110100000000" AFTER 25400 ns,
					"00000000000000000000000000000000" AFTER 25420 ns,
					"00000000000000000000110110000000" AFTER 25440 ns,
					"00000000000000000000000000000000" AFTER 25460 ns,
					"00000000000000000000111000000000" AFTER 25480 ns,
					"00000000000000000000000000000000" AFTER 25500 ns,
					"00000000000000000000111010000000" AFTER 25520 ns,
					"00000000000000000000000000000000" AFTER 25540 ns,
					"00000000000000000000111100000000" AFTER 25560 ns,
					"00000000000000000000000000000000" AFTER 25580 ns,
					"00000000000000000000111110000000" AFTER 25600 ns,
					"00000000000000000000000000000000" AFTER 25620 ns,
					"00000000000000000000000000000000" AFTER 25640 ns,
					"00000000000000000000000000000000" AFTER 25660 ns,
					"00000000000000001000000000000000" AFTER 25680 ns,
					"00000000000000000000000000000000" AFTER 25700 ns,
					"00000000000000010000000000000000" AFTER 25720 ns,
					"00000000000000000000000000000000" AFTER 25740 ns,
					"00000000000000011000000000000000" AFTER 25760 ns,
					"00000000000000000000000000000000" AFTER 25780 ns,
					"00000000000000100000000000000000" AFTER 25800 ns,
					"00000000000000000000000000000000" AFTER 25820 ns,
					"00000000000000101000000000000000" AFTER 25840 ns,
					"00000000000000000000000000000000" AFTER 25860 ns,
					"00000000000000110000000000000000" AFTER 25880 ns,
					"00000000000000000000000000000000" AFTER 25900 ns,
					"00000000000000111000000000000000" AFTER 25920 ns,
					"00000000000000000000000000000000" AFTER 25940 ns,
					"00000000000001000000000000000000" AFTER 25960 ns,
					"00000000000000000000000000000000" AFTER 25980 ns,
					"00000000000001001000000000000000" AFTER 26000 ns,
					"00000000000000000000000000000000" AFTER 26020 ns,
					"00000000000001010000000000000000" AFTER 26040 ns,
					"00000000000000000000000000000000" AFTER 26060 ns,
					"00000000000001011000000000000000" AFTER 26080 ns,
					"00000000000000000000000000000000" AFTER 26100 ns,
					"00000000000001100000000000000000" AFTER 26120 ns,
					"00000000000000000000000000000000" AFTER 26140 ns,
					"00000000000001101000000000000000" AFTER 26160 ns,
					"00000000000000000000000000000000" AFTER 26180 ns,
					"00000000000001110000000000000000" AFTER 26200 ns,
					"00000000000000000000000000000000" AFTER 26220 ns,
					"00000000000001111000000000000000" AFTER 26240 ns,
					"00000000000000000000000000000000" AFTER 26260 ns,
					"00000000000010000000000000000000" AFTER 26280 ns,
					"00000000000000000000000000000000" AFTER 26300 ns,
					"00000000000010001000000000000000" AFTER 26320 ns,
					"00000000000000000000000000000000" AFTER 26340 ns,
					"00000000000010010000000000000000" AFTER 26360 ns,
					"00000000000000000000000000000000" AFTER 26380 ns,
					"00000000000010011000000000000000" AFTER 26400 ns,
					"00000000000000000000000000000000" AFTER 26420 ns,
					"00000000000010100000000000000000" AFTER 26440 ns,
					"00000000000000000000000000000000" AFTER 26460 ns,
					"00000000000010101000000000000000" AFTER 26480 ns,
					"00000000000000000000000000000000" AFTER 26500 ns,
					"00000000000010110000000000000000" AFTER 26520 ns,
					"00000000000000000000000000000000" AFTER 26540 ns,
					"00000000000010111000000000000000" AFTER 26560 ns,
					"00000000000000000000000000000000" AFTER 26580 ns,
					"00000000000011000000000000000000" AFTER 26600 ns,
					"00000000000000000000000000000000" AFTER 26620 ns,
					"00000000000011001000000000000000" AFTER 26640 ns,
					"00000000000000000000000000000000" AFTER 26660 ns,
					"00000000000011010000000000000000" AFTER 26680 ns,
					"00000000000000000000000000000000" AFTER 26700 ns,
					"00000000000011011000000000000000" AFTER 26720 ns,
					"00000000000000000000000000000000" AFTER 26740 ns,
					"00000000000011100000000000000000" AFTER 26760 ns,
					"00000000000000000000000000000000" AFTER 26780 ns,
					"00000000000011101000000000000000" AFTER 26800 ns,
					"00000000000000000000000000000000" AFTER 26820 ns,
					"00000000000011110000000000000000" AFTER 26840 ns,
					"00000000000000000000000000000000" AFTER 26860 ns,
					"00000000000011111000000000000000" AFTER 26880 ns,
					"00000000000000000000000000000000" AFTER 26900 ns,
					"00000000000000000000000000000000" AFTER 26920 ns,
					"00000000000000000000000000000000" AFTER 26940 ns,
					"00000000000000000000000010000000" AFTER 26960 ns,
					"00000000000000000000000000000000" AFTER 26980 ns,
					"00000000000000000000000100000000" AFTER 27000 ns,
					"00000000000000000000000000000000" AFTER 27020 ns,
					"00000000000000000000000110000000" AFTER 27040 ns,
					"00000000000000000000000000000000" AFTER 27060 ns,
					"00000000000000000000001000000000" AFTER 27080 ns,
					"00000000000000000000000000000000" AFTER 27100 ns,
					"00000000000000000000001010000000" AFTER 27120 ns,
					"00000000000000000000000000000000" AFTER 27140 ns,
					"00000000000000000000001100000000" AFTER 27160 ns,
					"00000000000000000000000000000000" AFTER 27180 ns,
					"00000000000000000000001110000000" AFTER 27200 ns,
					"00000000000000000000000000000000" AFTER 27220 ns,
					"00000000000000000000010000000000" AFTER 27240 ns,
					"00000000000000000000000000000000" AFTER 27260 ns,
					"00000000000000000000010010000000" AFTER 27280 ns,
					"00000000000000000000000000000000" AFTER 27300 ns,
					"00000000000000000000010100000000" AFTER 27320 ns,
					"00000000000000000000000000000000" AFTER 27340 ns,
					"00000000000000000000010110000000" AFTER 27360 ns,
					"00000000000000000000000000000000" AFTER 27380 ns,
					"00000000000000000000011000000000" AFTER 27400 ns,
					"00000000000000000000000000000000" AFTER 27420 ns,
					"00000000000000000000011010000000" AFTER 27440 ns,
					"00000000000000000000000000000000" AFTER 27460 ns,
					"00000000000000000000011100000000" AFTER 27480 ns,
					"00000000000000000000000000000000" AFTER 27500 ns,
					"00000000000000000000011110000000" AFTER 27520 ns,
					"00000000000000000000000000000000" AFTER 27540 ns,
					"00000000000000000000100000000000" AFTER 27560 ns,
					"00000000000000000000000000000000" AFTER 27580 ns,
					"00000000000000000000100010000000" AFTER 27600 ns,
					"00000000000000000000000000000000" AFTER 27620 ns,
					"00000000000000000000100100000000" AFTER 27640 ns,
					"00000000000000000000000000000000" AFTER 27660 ns,
					"00000000000000000000100110000000" AFTER 27680 ns,
					"00000000000000000000000000000000" AFTER 27700 ns,
					"00000000000000000000101000000000" AFTER 27720 ns,
					"00000000000000000000000000000000" AFTER 27740 ns,
					"00000000000000000000101010000000" AFTER 27760 ns,
					"00000000000000000000000000000000" AFTER 27780 ns,
					"00000000000000000000101100000000" AFTER 27800 ns,
					"00000000000000000000000000000000" AFTER 27820 ns,
					"00000000000000000000101110000000" AFTER 27840 ns,
					"00000000000000000000000000000000" AFTER 27860 ns,
					"00000000000000000000110000000000" AFTER 27880 ns,
					"00000000000000000000000000000000" AFTER 27900 ns,
					"00000000000000000000110010000000" AFTER 27920 ns,
					"00000000000000000000000000000000" AFTER 27940 ns,
					"00000000000000000000110100000000" AFTER 27960 ns,
					"00000000000000000000000000000000" AFTER 27980 ns,
					"00000000000000000000110110000000" AFTER 28000 ns,
					"00000000000000000000000000000000" AFTER 28020 ns,
					"00000000000000000000111000000000" AFTER 28040 ns,
					"00000000000000000000000000000000" AFTER 28060 ns,
					"00000000000000000000111010000000" AFTER 28080 ns,
					"00000000000000000000000000000000" AFTER 28100 ns,
					"00000000000000000000111100000000" AFTER 28120 ns,
					"00000000000000000000000000000000" AFTER 28140 ns,
					"00000000000000000000111110000000" AFTER 28160 ns,
					"00000000000000000000000000000000" AFTER 28180 ns,
					"00000000000000000000000000000000" AFTER 28200 ns,
					"00000000000000000000000000000000" AFTER 28220 ns,
					"00000000000000000000000000000000" AFTER 28240 ns,
					"00000000000000000000000000000000" AFTER 28260 ns,
					"00000000000000000000000000000000" AFTER 28280 ns,
					"00000000000000000000000000000000" AFTER 28300 ns,
					"00000000000000000000000000000000" AFTER 28320 ns,
					"00000000000000000000000000000000" AFTER 28340 ns,
					"00000000000000000000000000000000" AFTER 28360 ns,
					"00000000000000000000000000000000" AFTER 28380 ns,
					"00000000000000000000000000000100" AFTER 28400 ns,
					"00000000000000000000000000000000" AFTER 28420 ns,
					"00000000000000000000000000001000" AFTER 28440 ns,
					"00000000000000000000000000000000" AFTER 28460 ns,
					"00000000000000000000000000001100" AFTER 28480 ns,
					"00000000000000000000000000000000" AFTER 28500 ns,
					"00000000000000000000000000010000" AFTER 28520 ns,
					"00000000000000000000000000000000" AFTER 28540 ns,
					"00000000000000000000000000010100" AFTER 28560 ns,
					"00000000000000000000000000000000" AFTER 28580 ns,
					"00000000000000000000000000011000" AFTER 28600 ns,
					"00000000000000000000000000000000" AFTER 28620 ns,
					"00000000000000000000000000011100" AFTER 28640 ns,
					"00000000000000000000000000000000" AFTER 28660 ns,
					"00000000000000000000000000100000" AFTER 28680 ns,
					"00000000000000000000000000000000" AFTER 28700 ns,
					"00000000000000000000000000100100" AFTER 28720 ns,
					"00000000000000000000000000000000" AFTER 28740 ns,
					"00000000000000000000000000101000" AFTER 28760 ns,
					"00000000000000000000000000000000" AFTER 28780 ns,
					"00000000000000000000000000101100" AFTER 28800 ns,
					"00000000000000000000000000000000" AFTER 28820 ns,
					"00000000000000000000000000110000" AFTER 28840 ns,
					"00000000000000000000000000000000" AFTER 28860 ns,
					"00000000000000000000000000110100" AFTER 28880 ns,
					"00000000000000000000000000000000" AFTER 28900 ns,
					"00000000000000000000000000111000" AFTER 28920 ns,
					"00000000000000000000000000000000" AFTER 28940 ns,
					"00000000000000000000000000111100" AFTER 28960 ns,
					"00000000000000000000000000000000" AFTER 28980 ns,
					"00000000000000000000000001000000" AFTER 29000 ns,
					"00000000000000000000000000000000" AFTER 29020 ns,
					"00000000000000000000000001000100" AFTER 29040 ns,
					"00000000000000000000000000000000" AFTER 29060 ns,
					"00000000000000000000000001001000" AFTER 29080 ns,
					"00000000000000000000000000000000" AFTER 29100 ns,
					"00000000000000000000000001001100" AFTER 29120 ns,
					"00000000000000000000000000000000" AFTER 29140 ns,
					"00000000000000000000000001010000" AFTER 29160 ns,
					"00000000000000000000000000000000" AFTER 29180 ns,
					"00000000000000000000000001010100" AFTER 29200 ns,
					"00000000000000000000000000000000" AFTER 29220 ns,
					"00000000000000000000000001011000" AFTER 29240 ns,
					"00000000000000000000000000000000" AFTER 29260 ns,
					"00000000000000000000000001011100" AFTER 29280 ns,
					"00000000000000000000000000000000" AFTER 29300 ns,
					"00000000000000000000000001100000" AFTER 29320 ns,
					"00000000000000000000000000000000" AFTER 29340 ns,
					"00000000000000000000000001100100" AFTER 29360 ns,
					"00000000000000000000000000000000" AFTER 29380 ns,
					"00000000000000000000000001101000" AFTER 29400 ns,
					"00000000000000000000000000000000" AFTER 29420 ns,
					"00000000000000000000000001101100" AFTER 29440 ns,
					"00000000000000000000000000000000" AFTER 29460 ns,
					"00000000000000000000000001110000" AFTER 29480 ns,
					"00000000000000000000000000000000" AFTER 29500 ns,
					"00000000000000000000000001110100" AFTER 29520 ns,
					"00000000000000000000000000000000" AFTER 29540 ns,
					"00000000000000000000000001111000" AFTER 29560 ns,
					"00000000000000000000000000000000" AFTER 29580 ns,
					"00000000000000000000000001111100" AFTER 29600 ns,
					"00000000000000000000000000000000" AFTER 29620 ns,
					"00000000000000000000000000000000" AFTER 29640 ns,
					"00000000000000000000000000000000" AFTER 29660 ns,
					"00000000000000000000000000000000" AFTER 29680 ns,
					"00000000000000000000000000000000" AFTER 29700 ns,
					"00000000000100000000000000000000" AFTER 29720 ns,
					"00000000000000000000000000000000" AFTER 29740 ns,
					"00000000001000000000000000000000" AFTER 29760 ns,
					"00000000000000000000000000000000" AFTER 29780 ns,
					"00000000001100000000000000000000" AFTER 29800 ns,
					"00000000000000000000000000000000" AFTER 29820 ns,
					"00000000010000000000000000000000" AFTER 29840 ns,
					"00000000000000000000000000000000" AFTER 29860 ns,
					"00000000010100000000000000000000" AFTER 29880 ns,
					"00000000000000000000000000000000" AFTER 29900 ns,
					"00000000011000000000000000000000" AFTER 29920 ns,
					"00000000000000000000000000000000" AFTER 29940 ns,
					"00000000011100000000000000000000" AFTER 29960 ns,
					"00000000000000000000000000000000" AFTER 29980 ns,
					"00000000100000000000000000000000" AFTER 30000 ns,
					"00000000000000000000000000000000" AFTER 30020 ns,
					"00000000100100000000000000000000" AFTER 30040 ns,
					"00000000000000000000000000000000" AFTER 30060 ns,
					"00000000101000000000000000000000" AFTER 30080 ns,
					"00000000000000000000000000000000" AFTER 30100 ns,
					"00000000101100000000000000000000" AFTER 30120 ns,
					"00000000000000000000000000000000" AFTER 30140 ns,
					"00000000110000000000000000000000" AFTER 30160 ns,
					"00000000000000000000000000000000" AFTER 30180 ns,
					"00000000110100000000000000000000" AFTER 30200 ns,
					"00000000000000000000000000000000" AFTER 30220 ns,
					"00000000111000000000000000000000" AFTER 30240 ns,
					"00000000000000000000000000000000" AFTER 30260 ns,
					"00000000111100000000000000000000" AFTER 30280 ns,
					"00000000000000000000000000000000" AFTER 30300 ns,
					"00000001000000000000000000000000" AFTER 30320 ns,
					"00000000000000000000000000000000" AFTER 30340 ns,
					"00000001000100000000000000000000" AFTER 30360 ns,
					"00000000000000000000000000000000" AFTER 30380 ns,
					"00000001001000000000000000000000" AFTER 30400 ns,
					"00000000000000000000000000000000" AFTER 30420 ns,
					"00000001001100000000000000000000" AFTER 30440 ns,
					"00000000000000000000000000000000" AFTER 30460 ns,
					"00000001010000000000000000000000" AFTER 30480 ns,
					"00000000000000000000000000000000" AFTER 30500 ns,
					"00000001010100000000000000000000" AFTER 30520 ns,
					"00000000000000000000000000000000" AFTER 30540 ns,
					"00000001011000000000000000000000" AFTER 30560 ns,
					"00000000000000000000000000000000" AFTER 30580 ns,
					"00000001011100000000000000000000" AFTER 30600 ns,
					"00000000000000000000000000000000" AFTER 30620 ns,
					"00000001100000000000000000000000" AFTER 30640 ns,
					"00000000000000000000000000000000" AFTER 30660 ns,
					"00000001100100000000000000000000" AFTER 30680 ns,
					"00000000000000000000000000000000" AFTER 30700 ns,
					"00000001101000000000000000000000" AFTER 30720 ns,
					"00000000000000000000000000000000" AFTER 30740 ns,
					"00000001101100000000000000000000" AFTER 30760 ns,
					"00000000000000000000000000000000" AFTER 30780 ns,
					"00000001110000000000000000000000" AFTER 30800 ns,
					"00000000000000000000000000000000" AFTER 30820 ns,
					"00000001110100000000000000000000" AFTER 30840 ns,
					"00000000000000000000000000000000" AFTER 30860 ns,
					"00000001111000000000000000000000" AFTER 30880 ns,
					"00000000000000000000000000000000" AFTER 30900 ns,
					"00000001111100000000000000000000" AFTER 30920 ns,
					"00000000000000000000000000000000" AFTER 30940 ns,
					"00000000000000000000000000000000" AFTER 30960 ns;

CsrRegisters <= x"00000000" AFTER 00020 ns,
x"00000533" AFTER 00040 ns,
x"00000000" AFTER 00060 ns,
x"0000052F" AFTER 00080 ns,
x"00000000" AFTER 00100 ns,
x"0000052B" AFTER 00120 ns,
x"00000000" AFTER 00140 ns,
x"00000527" AFTER 00160 ns,
x"00000000" AFTER 00180 ns,
x"00000523" AFTER 00200 ns,
x"00000000" AFTER 00220 ns,
x"0000051F" AFTER 00240 ns,
x"00000000" AFTER 00260 ns,
x"0000051B" AFTER 00280 ns,
x"00000000" AFTER 00300 ns,
x"00000517" AFTER 00320 ns,
x"00000000" AFTER 00340 ns,
x"00000513" AFTER 00360 ns,
x"00000000" AFTER 00380 ns,
x"0000050F" AFTER 00400 ns,
x"00000000" AFTER 00420 ns,
x"0000050B" AFTER 00440 ns,
x"00000000" AFTER 00460 ns,
x"00000507" AFTER 00480 ns,
x"00000000" AFTER 00500 ns,
x"00000503" AFTER 00520 ns,
x"00000000" AFTER 00540 ns,
x"000004FF" AFTER 00560 ns,
x"00000000" AFTER 00580 ns,
x"000004FB" AFTER 00600 ns,
x"00000000" AFTER 00620 ns,
x"000004F7" AFTER 00640 ns,
x"00000000" AFTER 00660 ns,
x"000004F3" AFTER 00680 ns,
x"00000000" AFTER 00700 ns,
x"000004EF" AFTER 00720 ns,
x"00000000" AFTER 00740 ns,
x"000004EB" AFTER 00760 ns,
x"00000000" AFTER 00780 ns,
x"000004E7" AFTER 00800 ns,
x"00000000" AFTER 00820 ns,
x"000004E3" AFTER 00840 ns,
x"00000000" AFTER 00860 ns,
x"000004DF" AFTER 00880 ns,
x"00000000" AFTER 00900 ns,
x"000004DB" AFTER 00920 ns,
x"00000000" AFTER 00940 ns,
x"000004D7" AFTER 00960 ns,
x"00000000" AFTER 00980 ns,
x"000004D3" AFTER 01000 ns,
x"00000000" AFTER 01020 ns,
x"000004CF" AFTER 01040 ns,
x"00000000" AFTER 01060 ns,
x"000004CB" AFTER 01080 ns,
x"00000000" AFTER 01100 ns,
x"000004C7" AFTER 01120 ns,
x"00000000" AFTER 01140 ns,
x"000004C3" AFTER 01160 ns,
x"00000000" AFTER 01180 ns,
x"000004BF" AFTER 01200 ns,
x"00000000" AFTER 01220 ns,
x"000004BB" AFTER 01240 ns,
x"00000000" AFTER 01260 ns,
x"000004B7" AFTER 01280 ns,
x"00000000" AFTER 01300 ns,
x"000004B3" AFTER 01320 ns,
x"00000000" AFTER 01340 ns,
x"000004AF" AFTER 01360 ns,
x"00000000" AFTER 01380 ns,
x"000004AB" AFTER 01400 ns,
x"00000000" AFTER 01420 ns,
x"000004A7" AFTER 01440 ns,
x"00000000" AFTER 01460 ns,
x"000004A3" AFTER 01480 ns,
x"00000000" AFTER 01500 ns,
x"0000049F" AFTER 01520 ns,
x"00000000" AFTER 01540 ns,
x"0000049B" AFTER 01560 ns,
x"00000000" AFTER 01580 ns,
x"00000497" AFTER 01600 ns,
x"00000000" AFTER 01620 ns,
x"00000493" AFTER 01640 ns,
x"00000000" AFTER 01660 ns,
x"0000048F" AFTER 01680 ns,
x"00000000" AFTER 01700 ns,
x"0000048B" AFTER 01720 ns,
x"00000000" AFTER 01740 ns,
x"00000487" AFTER 01760 ns,
x"00000000" AFTER 01780 ns,
x"00000483" AFTER 01800 ns,
x"00000000" AFTER 01820 ns,
x"0000047F" AFTER 01840 ns,
x"00000000" AFTER 01860 ns,
x"0000047B" AFTER 01880 ns,
x"00000000" AFTER 01900 ns,
x"00000477" AFTER 01920 ns,
x"00000000" AFTER 01940 ns,
x"00000473" AFTER 01960 ns,
x"00000000" AFTER 01980 ns,
x"0000046F" AFTER 02000 ns,
x"00000000" AFTER 02020 ns,
x"0000046B" AFTER 02040 ns,
x"00000000" AFTER 02060 ns,
x"00000467" AFTER 02080 ns,
x"00000000" AFTER 02100 ns,
x"00000463" AFTER 02120 ns,
x"00000000" AFTER 02140 ns,
x"0000045F" AFTER 02160 ns,
x"00000000" AFTER 02180 ns,
x"0000045B" AFTER 02200 ns,
x"00000000" AFTER 02220 ns,
x"00000457" AFTER 02240 ns,
x"00000000" AFTER 02260 ns,
x"00000453" AFTER 02280 ns,
x"00000000" AFTER 02300 ns,
x"0000044F" AFTER 02320 ns,
x"00000000" AFTER 02340 ns,
x"0000044B" AFTER 02360 ns,
x"00000000" AFTER 02380 ns,
x"00000447" AFTER 02400 ns,
x"00000000" AFTER 02420 ns,
x"00000443" AFTER 02440 ns,
x"00000000" AFTER 02460 ns,
x"0000043F" AFTER 02480 ns,
x"00000000" AFTER 02500 ns,
x"0000043B" AFTER 02520 ns,
x"00000000" AFTER 02540 ns,
x"00000437" AFTER 02560 ns,
x"00000000" AFTER 02580 ns,
x"00000433" AFTER 02600 ns,
x"00000000" AFTER 02620 ns,
x"0000042F" AFTER 02640 ns,
x"00000000" AFTER 02660 ns,
x"0000042B" AFTER 02680 ns,
x"00000000" AFTER 02700 ns,
x"00000427" AFTER 02720 ns,
x"00000000" AFTER 02740 ns,
x"00000423" AFTER 02760 ns,
x"00000000" AFTER 02780 ns,
x"0000041F" AFTER 02800 ns,
x"00000000" AFTER 02820 ns,
x"0000041B" AFTER 02840 ns,
x"00000000" AFTER 02860 ns,
x"00000417" AFTER 02880 ns,
x"00000000" AFTER 02900 ns,
x"00000413" AFTER 02920 ns,
x"00000000" AFTER 02940 ns,
x"0000040F" AFTER 02960 ns,
x"00000000" AFTER 02980 ns,
x"0000040B" AFTER 03000 ns,
x"00000000" AFTER 03020 ns,
x"00000407" AFTER 03040 ns,
x"00000000" AFTER 03060 ns,
x"00000403" AFTER 03080 ns,
x"00000000" AFTER 03100 ns,
x"000003FF" AFTER 03120 ns,
x"00000000" AFTER 03140 ns,
x"000003FB" AFTER 03160 ns,
x"00000000" AFTER 03180 ns,
x"000003F7" AFTER 03200 ns,
x"00000000" AFTER 03220 ns,
x"000003F3" AFTER 03240 ns,
x"00000000" AFTER 03260 ns,
x"000003EF" AFTER 03280 ns,
x"00000000" AFTER 03300 ns,
x"000003EB" AFTER 03320 ns,
x"00000000" AFTER 03340 ns,
x"000003E7" AFTER 03360 ns,
x"00000000" AFTER 03380 ns,
x"000003E3" AFTER 03400 ns,
x"00000000" AFTER 03420 ns,
x"000003DF" AFTER 03440 ns,
x"00000000" AFTER 03460 ns,
x"000003DB" AFTER 03480 ns,
x"00000000" AFTER 03500 ns,
x"000003D7" AFTER 03520 ns,
x"00000000" AFTER 03540 ns,
x"000003D3" AFTER 03560 ns,
x"00000000" AFTER 03580 ns,
x"000003CF" AFTER 03600 ns,
x"00000000" AFTER 03620 ns,
x"000003CB" AFTER 03640 ns,
x"00000000" AFTER 03660 ns,
x"000003C7" AFTER 03680 ns,
x"00000000" AFTER 03700 ns,
x"000003C3" AFTER 03720 ns,
x"00000000" AFTER 03740 ns,
x"000003BF" AFTER 03760 ns,
x"00000000" AFTER 03780 ns,
x"000003BB" AFTER 03800 ns,
x"00000000" AFTER 03820 ns,
x"000003B7" AFTER 03840 ns,
x"00000000" AFTER 03860 ns,
x"000003B3" AFTER 03880 ns,
x"00000000" AFTER 03900 ns,
x"000003AF" AFTER 03920 ns,
x"00000000" AFTER 03940 ns,
x"000003AB" AFTER 03960 ns,
x"00000000" AFTER 03980 ns,
x"000003A7" AFTER 04000 ns,
x"00000000" AFTER 04020 ns,
x"000003A3" AFTER 04040 ns,
x"00000000" AFTER 04060 ns,
x"0000039F" AFTER 04080 ns,
x"00000000" AFTER 04100 ns,
x"0000039B" AFTER 04120 ns,
x"00000000" AFTER 04140 ns,
x"00000397" AFTER 04160 ns,
x"00000000" AFTER 04180 ns,
x"00000393" AFTER 04200 ns,
x"00000000" AFTER 04220 ns,
x"0000038F" AFTER 04240 ns,
x"00000000" AFTER 04260 ns,
x"0000038B" AFTER 04280 ns,
x"00000000" AFTER 04300 ns,
x"00000387" AFTER 04320 ns,
x"00000000" AFTER 04340 ns,
x"00000383" AFTER 04360 ns,
x"00000000" AFTER 04380 ns,
x"0000037F" AFTER 04400 ns,
x"00000000" AFTER 04420 ns,
x"0000037B" AFTER 04440 ns,
x"00000000" AFTER 04460 ns,
x"00000377" AFTER 04480 ns,
x"00000000" AFTER 04500 ns,
x"00000373" AFTER 04520 ns,
x"00000000" AFTER 04540 ns,
x"0000036F" AFTER 04560 ns,
x"00000000" AFTER 04580 ns,
x"0000036B" AFTER 04600 ns,
x"00000000" AFTER 04620 ns,
x"00000367" AFTER 04640 ns,
x"00000000" AFTER 04660 ns,
x"00000363" AFTER 04680 ns,
x"00000000" AFTER 04700 ns,
x"0000035F" AFTER 04720 ns,
x"00000000" AFTER 04740 ns,
x"0000035B" AFTER 04760 ns,
x"00000000" AFTER 04780 ns,
x"00000357" AFTER 04800 ns,
x"00000000" AFTER 04820 ns,
x"00000353" AFTER 04840 ns,
x"00000000" AFTER 04860 ns,
x"0000034F" AFTER 04880 ns,
x"00000000" AFTER 04900 ns,
x"0000034B" AFTER 04920 ns,
x"00000000" AFTER 04940 ns,
x"00000347" AFTER 04960 ns,
x"00000000" AFTER 04980 ns,
x"00000343" AFTER 05000 ns,
x"00000000" AFTER 05020 ns,
x"0000033F" AFTER 05040 ns,
x"00000000" AFTER 05060 ns,
x"0000033B" AFTER 05080 ns,
x"00000000" AFTER 05100 ns,
x"00000337" AFTER 05120 ns,
x"00000000" AFTER 05140 ns,
x"00000333" AFTER 05160 ns,
x"00000000" AFTER 05180 ns,
x"0000032F" AFTER 05200 ns,
x"00000000" AFTER 05220 ns,
x"0000032B" AFTER 05240 ns,
x"00000000" AFTER 05260 ns,
x"00000327" AFTER 05280 ns,
x"00000000" AFTER 05300 ns,
x"00000323" AFTER 05320 ns,
x"00000000" AFTER 05340 ns,
x"0000031F" AFTER 05360 ns,
x"00000000" AFTER 05380 ns,
x"0000031B" AFTER 05400 ns,
x"00000000" AFTER 05420 ns,
x"00000317" AFTER 05440 ns,
x"00000000" AFTER 05460 ns,
x"00000313" AFTER 05480 ns,
x"00000000" AFTER 05500 ns,
x"0000030F" AFTER 05520 ns,
x"00000000" AFTER 05540 ns,
x"0000030B" AFTER 05560 ns,
x"00000000" AFTER 05580 ns,
x"00000307" AFTER 05600 ns,
x"00000000" AFTER 05620 ns,
x"00000303" AFTER 05640 ns,
x"00000000" AFTER 05660 ns,
x"000002FF" AFTER 05680 ns,
x"00000000" AFTER 05700 ns,
x"000002FB" AFTER 05720 ns,
x"00000000" AFTER 05740 ns,
x"000002F7" AFTER 05760 ns,
x"00000000" AFTER 05780 ns,
x"000002F3" AFTER 05800 ns,
x"00000000" AFTER 05820 ns,
x"000002EF" AFTER 05840 ns,
x"00000000" AFTER 05860 ns,
x"000002EB" AFTER 05880 ns,
x"00000000" AFTER 05900 ns,
x"000002E7" AFTER 05920 ns,
x"00000000" AFTER 05940 ns,
x"000002E3" AFTER 05960 ns,
x"00000000" AFTER 05980 ns,
x"000002DF" AFTER 06000 ns,
x"00000000" AFTER 06020 ns,
x"000002DB" AFTER 06040 ns,
x"00000000" AFTER 06060 ns,
x"000002D7" AFTER 06080 ns,
x"00000000" AFTER 06100 ns,
x"000002D3" AFTER 06120 ns,
x"00000000" AFTER 06140 ns,
x"000002CF" AFTER 06160 ns,
x"00000000" AFTER 06180 ns,
x"000002CB" AFTER 06200 ns,
x"00000000" AFTER 06220 ns,
x"000002C7" AFTER 06240 ns,
x"00000000" AFTER 06260 ns,
x"000002C3" AFTER 06280 ns,
x"00000000" AFTER 06300 ns,
x"000002BF" AFTER 06320 ns,
x"00000000" AFTER 06340 ns,
x"000002BB" AFTER 06360 ns,
x"00000000" AFTER 06380 ns,
x"000002B7" AFTER 06400 ns,
x"00000000" AFTER 06420 ns,
x"000002B3" AFTER 06440 ns,
x"00000000" AFTER 06460 ns,
x"000002AF" AFTER 06480 ns,
x"00000000" AFTER 06500 ns,
x"000002AB" AFTER 06520 ns,
x"00000000" AFTER 06540 ns,
x"000002A7" AFTER 06560 ns,
x"00000000" AFTER 06580 ns,
x"000002A3" AFTER 06600 ns,
x"00000000" AFTER 06620 ns,
x"0000029F" AFTER 06640 ns,
x"00000000" AFTER 06660 ns,
x"0000029B" AFTER 06680 ns,
x"00000000" AFTER 06700 ns,
x"00000297" AFTER 06720 ns,
x"00000000" AFTER 06740 ns,
x"00000293" AFTER 06760 ns,
x"00000000" AFTER 06780 ns,
x"0000028F" AFTER 06800 ns,
x"00000000" AFTER 06820 ns,
x"0000028B" AFTER 06840 ns,
x"00000000" AFTER 06860 ns,
x"00000287" AFTER 06880 ns,
x"00000000" AFTER 06900 ns,
x"00000283" AFTER 06920 ns,
x"00000000" AFTER 06940 ns,
x"0000027F" AFTER 06960 ns,
x"00000000" AFTER 06980 ns,
x"0000027B" AFTER 07000 ns,
x"00000000" AFTER 07020 ns,
x"00000277" AFTER 07040 ns,
x"00000000" AFTER 07060 ns,
x"00000273" AFTER 07080 ns,
x"00000000" AFTER 07100 ns,
x"0000026F" AFTER 07120 ns,
x"00000000" AFTER 07140 ns,
x"0000026B" AFTER 07160 ns,
x"00000000" AFTER 07180 ns,
x"00000267" AFTER 07200 ns,
x"00000000" AFTER 07220 ns,
x"00000263" AFTER 07240 ns,
x"00000000" AFTER 07260 ns,
x"0000025F" AFTER 07280 ns,
x"00000000" AFTER 07300 ns,
x"0000025B" AFTER 07320 ns,
x"00000000" AFTER 07340 ns,
x"00000257" AFTER 07360 ns,
x"00000000" AFTER 07380 ns,
x"00000253" AFTER 07400 ns,
x"00000000" AFTER 07420 ns,
x"0000024F" AFTER 07440 ns,
x"00000000" AFTER 07460 ns,
x"0000024B" AFTER 07480 ns,
x"00000000" AFTER 07500 ns,
x"00000247" AFTER 07520 ns,
x"00000000" AFTER 07540 ns,
x"00000243" AFTER 07560 ns,
x"00000000" AFTER 07580 ns,
x"0000023F" AFTER 07600 ns,
x"00000000" AFTER 07620 ns,
x"0000023B" AFTER 07640 ns,
x"00000000" AFTER 07660 ns,
x"00000237" AFTER 07680 ns,
x"00000000" AFTER 07700 ns,
x"00000233" AFTER 07720 ns,
x"00000000" AFTER 07740 ns,
x"0000022F" AFTER 07760 ns,
x"00000000" AFTER 07780 ns,
x"0000022B" AFTER 07800 ns,
x"00000000" AFTER 07820 ns,
x"00000227" AFTER 07840 ns,
x"00000000" AFTER 07860 ns,
x"00000223" AFTER 07880 ns,
x"00000000" AFTER 07900 ns,
x"0000021F" AFTER 07920 ns,
x"00000000" AFTER 07940 ns,
x"0000021B" AFTER 07960 ns,
x"00000000" AFTER 07980 ns,
x"00000217" AFTER 08000 ns,
x"00000000" AFTER 08020 ns,
x"00000213" AFTER 08040 ns,
x"00000000" AFTER 08060 ns,
x"0000020F" AFTER 08080 ns,
x"00000000" AFTER 08100 ns,
x"0000020B" AFTER 08120 ns,
x"00000000" AFTER 08140 ns,
x"00000207" AFTER 08160 ns,
x"00000000" AFTER 08180 ns,
x"00000203" AFTER 08200 ns,
x"00000000" AFTER 08220 ns,
x"000001FF" AFTER 08240 ns,
x"00000000" AFTER 08260 ns,
x"000001FB" AFTER 08280 ns,
x"00000000" AFTER 08300 ns,
x"000001F7" AFTER 08320 ns,
x"00000000" AFTER 08340 ns,
x"000001F3" AFTER 08360 ns,
x"00000000" AFTER 08380 ns,
x"000001EF" AFTER 08400 ns,
x"00000000" AFTER 08420 ns,
x"000001EB" AFTER 08440 ns,
x"00000000" AFTER 08460 ns,
x"000001E7" AFTER 08480 ns,
x"00000000" AFTER 08500 ns,
x"000001E3" AFTER 08520 ns,
x"00000000" AFTER 08540 ns,
x"000001DF" AFTER 08560 ns,
x"00000000" AFTER 08580 ns,
x"000001DB" AFTER 08600 ns,
x"00000000" AFTER 08620 ns,
x"000001D7" AFTER 08640 ns,
x"00000000" AFTER 08660 ns,
x"000001D3" AFTER 08680 ns,
x"00000000" AFTER 08700 ns,
x"000001CF" AFTER 08720 ns,
x"00000000" AFTER 08740 ns,
x"000001CB" AFTER 08760 ns,
x"00000000" AFTER 08780 ns,
x"000001C7" AFTER 08800 ns,
x"00000000" AFTER 08820 ns,
x"000001C3" AFTER 08840 ns,
x"00000000" AFTER 08860 ns,
x"000001BF" AFTER 08880 ns,
x"00000000" AFTER 08900 ns,
x"000001BB" AFTER 08920 ns,
x"00000000" AFTER 08940 ns,
x"000001B7" AFTER 08960 ns,
x"00000000" AFTER 08980 ns,
x"000001B3" AFTER 09000 ns,
x"00000000" AFTER 09020 ns,
x"000001AF" AFTER 09040 ns,
x"00000000" AFTER 09060 ns,
x"000001AB" AFTER 09080 ns,
x"00000000" AFTER 09100 ns,
x"000001A7" AFTER 09120 ns,
x"00000000" AFTER 09140 ns,
x"000001A3" AFTER 09160 ns,
x"00000000" AFTER 09180 ns,
x"0000019F" AFTER 09200 ns,
x"00000000" AFTER 09220 ns,
x"0000019B" AFTER 09240 ns,
x"00000000" AFTER 09260 ns,
x"00000197" AFTER 09280 ns,
x"00000000" AFTER 09300 ns,
x"00000193" AFTER 09320 ns,
x"00000000" AFTER 09340 ns,
x"0000018F" AFTER 09360 ns,
x"00000000" AFTER 09380 ns,
x"0000018B" AFTER 09400 ns,
x"00000000" AFTER 09420 ns,
x"00000187" AFTER 09440 ns,
x"00000000" AFTER 09460 ns,
x"00000183" AFTER 09480 ns,
x"00000000" AFTER 09500 ns,
x"0000017F" AFTER 09520 ns,
x"00000000" AFTER 09540 ns,
x"0000017B" AFTER 09560 ns,
x"00000000" AFTER 09580 ns,
x"00000177" AFTER 09600 ns,
x"00000000" AFTER 09620 ns,
x"00000173" AFTER 09640 ns,
x"00000000" AFTER 09660 ns,
x"0000016F" AFTER 09680 ns,
x"00000000" AFTER 09700 ns,
x"0000016B" AFTER 09720 ns,
x"00000000" AFTER 09740 ns,
x"00000167" AFTER 09760 ns,
x"00000000" AFTER 09780 ns,
x"00000163" AFTER 09800 ns,
x"00000000" AFTER 09820 ns,
x"0000015F" AFTER 09840 ns,
x"00000000" AFTER 09860 ns,
x"0000015B" AFTER 09880 ns,
x"00000000" AFTER 09900 ns,
x"00000157" AFTER 09920 ns,
x"00000000" AFTER 09940 ns,
x"00000153" AFTER 09960 ns,
x"00000000" AFTER 09980 ns,
x"0000014F" AFTER 10000 ns,
x"00000000" AFTER 10020 ns,
x"0000014B" AFTER 10040 ns,
x"00000000" AFTER 10060 ns,
x"00000147" AFTER 10080 ns,
x"00000000" AFTER 10100 ns,
x"00000143" AFTER 10120 ns,
x"00000000" AFTER 10140 ns,
x"0000013F" AFTER 10160 ns,
x"00000000" AFTER 10180 ns,
x"0000013B" AFTER 10200 ns,
x"00000000" AFTER 10220 ns,
x"00000137" AFTER 10240 ns,
x"00000000" AFTER 10260 ns,
x"00000133" AFTER 10280 ns,
x"00000000" AFTER 10300 ns,
x"0000012F" AFTER 10320 ns,
x"00000000" AFTER 10340 ns,
x"0000012B" AFTER 10360 ns,
x"00000000" AFTER 10380 ns,
x"00000127" AFTER 10400 ns,
x"00000000" AFTER 10420 ns,
x"00000123" AFTER 10440 ns,
x"00000000" AFTER 10460 ns,
x"0000011F" AFTER 10480 ns,
x"00000000" AFTER 10500 ns,
x"0000011B" AFTER 10520 ns,
x"00000000" AFTER 10540 ns,
x"00000117" AFTER 10560 ns,
x"00000000" AFTER 10580 ns,
x"00000113" AFTER 10600 ns,
x"00000000" AFTER 10620 ns,
x"0000010F" AFTER 10640 ns,
x"00000000" AFTER 10660 ns,
x"0000010B" AFTER 10680 ns,
x"00000000" AFTER 10700 ns,
x"00000107" AFTER 10720 ns,
x"00000000" AFTER 10740 ns,
x"00000103" AFTER 10760 ns,
x"00000000" AFTER 10780 ns,
x"000000FF" AFTER 10800 ns,
x"00000000" AFTER 10820 ns,
x"000000FB" AFTER 10840 ns,
x"00000000" AFTER 10860 ns,
x"000000F7" AFTER 10880 ns,
x"00000000" AFTER 10900 ns,
x"000000F3" AFTER 10920 ns,
x"00000000" AFTER 10940 ns,
x"000000EF" AFTER 10960 ns,
x"00000000" AFTER 10980 ns,
x"000000EB" AFTER 11000 ns,
x"00000000" AFTER 11020 ns,
x"000000E7" AFTER 11040 ns,
x"00000000" AFTER 11060 ns,
x"000000E3" AFTER 11080 ns,
x"00000000" AFTER 11100 ns,
x"000000DF" AFTER 11120 ns,
x"00000000" AFTER 11140 ns,
x"000000DB" AFTER 11160 ns,
x"00000000" AFTER 11180 ns,
x"000000D7" AFTER 11200 ns,
x"00000000" AFTER 11220 ns,
x"000000D3" AFTER 11240 ns,
x"00000000" AFTER 11260 ns,
x"000000CF" AFTER 11280 ns,
x"00000000" AFTER 11300 ns,
x"000000CB" AFTER 11320 ns,
x"00000000" AFTER 11340 ns,
x"000000C7" AFTER 11360 ns,
x"00000000" AFTER 11380 ns,
x"000000C3" AFTER 11400 ns,
x"00000000" AFTER 11420 ns,
x"000000BF" AFTER 11440 ns,
x"00000000" AFTER 11460 ns,
x"000000BB" AFTER 11480 ns,
x"00000000" AFTER 11500 ns,
x"000000B7" AFTER 11520 ns,
x"00000000" AFTER 11540 ns,
x"000000B3" AFTER 11560 ns,
x"00000000" AFTER 11580 ns,
x"000000AF" AFTER 11600 ns,
x"00000000" AFTER 11620 ns,
x"000000AB" AFTER 11640 ns,
x"00000000" AFTER 11660 ns,
x"000000A7" AFTER 11680 ns,
x"00000000" AFTER 11700 ns,
x"000000A3" AFTER 11720 ns,
x"00000000" AFTER 11740 ns,
x"0000009F" AFTER 11760 ns,
x"00000000" AFTER 11780 ns,
x"0000009B" AFTER 11800 ns,
x"00000000" AFTER 11820 ns,
x"00000097" AFTER 11840 ns,
x"00000000" AFTER 11860 ns,
x"00000093" AFTER 11880 ns,
x"00000000" AFTER 11900 ns,
x"0000008F" AFTER 11920 ns,
x"00000000" AFTER 11940 ns,
x"0000008B" AFTER 11960 ns,
x"00000000" AFTER 11980 ns,
x"00000087" AFTER 12000 ns,
x"00000000" AFTER 12020 ns,
x"00000083" AFTER 12040 ns,
x"00000000" AFTER 12060 ns,
x"0000007F" AFTER 12080 ns,
x"00000000" AFTER 12100 ns,
x"0000007B" AFTER 12120 ns,
x"00000000" AFTER 12140 ns,
x"00000077" AFTER 12160 ns,
x"00000000" AFTER 12180 ns,
x"00000073" AFTER 12200 ns,
x"00000000" AFTER 12220 ns,
x"0000006F" AFTER 12240 ns,
x"00000000" AFTER 12260 ns,
x"0000006B" AFTER 12280 ns,
x"00000000" AFTER 12300 ns,
x"00000067" AFTER 12320 ns,
x"00000000" AFTER 12340 ns,
x"00000063" AFTER 12360 ns,
x"00000000" AFTER 12380 ns,
x"0000005F" AFTER 12400 ns,
x"00000000" AFTER 12420 ns,
x"0000005B" AFTER 12440 ns,
x"00000000" AFTER 12460 ns,
x"00000057" AFTER 12480 ns,
x"00000000" AFTER 12500 ns,
x"00000053" AFTER 12520 ns,
x"00000000" AFTER 12540 ns,
x"0000004F" AFTER 12560 ns,
x"00000000" AFTER 12580 ns,
x"0000004B" AFTER 12600 ns,
x"00000000" AFTER 12620 ns,
x"00000047" AFTER 12640 ns,
x"00000000" AFTER 12660 ns,
x"00000043" AFTER 12680 ns,
x"00000000" AFTER 12700 ns,
x"0000003F" AFTER 12720 ns,
x"00000000" AFTER 12740 ns,
x"0000003B" AFTER 12760 ns,
x"00000000" AFTER 12780 ns,
x"00000037" AFTER 12800 ns,
x"00000000" AFTER 12820 ns,
x"00000033" AFTER 12840 ns,
x"00000000" AFTER 12860 ns,
x"0000002F" AFTER 12880 ns,
x"00000000" AFTER 12900 ns,
x"0000002B" AFTER 12920 ns,
x"00000000" AFTER 12940 ns,
x"00000027" AFTER 12960 ns,
x"00000000" AFTER 12980 ns,
x"00000023" AFTER 13000 ns,
x"00000000" AFTER 13020 ns,
x"0000001F" AFTER 13040 ns,
x"00000000" AFTER 13060 ns,
x"0000001B" AFTER 13080 ns,
x"00000000" AFTER 13100 ns,
x"00000017" AFTER 13120 ns,
x"00000000" AFTER 13140 ns,
x"00000013" AFTER 13160 ns,
x"00000000" AFTER 13180 ns,
x"0000000F" AFTER 13200 ns,
x"00000000" AFTER 13220 ns,
x"0000000B" AFTER 13240 ns,
x"00000000" AFTER 13260 ns,
x"00000007" AFTER 13280 ns,
x"00000000" AFTER 13300 ns,
x"00000003" AFTER 13320 ns,
x"00000000" AFTER 13340 ns,
x"EE6B27FB" AFTER 13360 ns,
x"00000000" AFTER 13380 ns,
x"EE6B27F7" AFTER 13400 ns,
x"00000000" AFTER 13420 ns,
x"EE6B27F3" AFTER 13440 ns,
x"00000000" AFTER 13460 ns,
x"EE6B27EF" AFTER 13480 ns,
x"00000000" AFTER 13500 ns,
x"EE6B27EB" AFTER 13520 ns,
x"00000000" AFTER 13540 ns,
x"EE6B27E7" AFTER 13560 ns,
x"00000000" AFTER 13580 ns,
x"EE6B27E3" AFTER 13600 ns,
x"00000000" AFTER 13620 ns,
x"EE6B27DF" AFTER 13640 ns,
x"00000000" AFTER 13660 ns,
x"EE6B27DB" AFTER 13680 ns,
x"00000000" AFTER 13700 ns,
x"EE6B27D7" AFTER 13720 ns,
x"00000000" AFTER 13740 ns,
x"EE6B27D3" AFTER 13760 ns,
x"00000000" AFTER 13780 ns,
x"EE6B27CF" AFTER 13800 ns,
x"00000000" AFTER 13820 ns,
x"EE6B27CB" AFTER 13840 ns,
x"00000000" AFTER 13860 ns,
x"EE6B27C7" AFTER 13880 ns,
x"00000000" AFTER 13900 ns,
x"EE6B27C3" AFTER 13920 ns,
x"00000000" AFTER 13940 ns,
x"EE6B27BF" AFTER 13960 ns,
x"00000000" AFTER 13980 ns,
x"EE6B27BB" AFTER 14000 ns,
x"00000000" AFTER 14020 ns,
x"EE6B27B7" AFTER 14040 ns,
x"00000000" AFTER 14060 ns,
x"EE6B27B3" AFTER 14080 ns,
x"00000000" AFTER 14100 ns,
x"EE6B27AF" AFTER 14120 ns,
x"00000000" AFTER 14140 ns,
x"EE6B27AB" AFTER 14160 ns,
x"00000000" AFTER 14180 ns,
x"EE6B27A7" AFTER 14200 ns,
x"00000000" AFTER 14220 ns,
x"EE6B27A3" AFTER 14240 ns,
x"00000000" AFTER 14260 ns,
x"EE6B279F" AFTER 14280 ns,
x"00000000" AFTER 14300 ns,
x"EE6B279B" AFTER 14320 ns,
x"00000000" AFTER 14340 ns,
x"EE6B2797" AFTER 14360 ns,
x"00000000" AFTER 14380 ns,
x"EE6B2793" AFTER 14400 ns,
x"00000000" AFTER 14420 ns,
x"EE6B278F" AFTER 14440 ns,
x"00000000" AFTER 14460 ns,
x"EE6B278B" AFTER 14480 ns,
x"00000000" AFTER 14500 ns,
x"EE6B2787" AFTER 14520 ns,
x"00000000" AFTER 14540 ns,
x"EE6B2783" AFTER 14560 ns,
x"00000000" AFTER 14580 ns,
x"EE6B277F" AFTER 14600 ns,
x"00000000" AFTER 14620 ns,
x"EE6B277B" AFTER 14640 ns,
x"00000000" AFTER 14660 ns,
x"EE6B2777" AFTER 14680 ns,
x"00000000" AFTER 14700 ns,
x"EE6B2773" AFTER 14720 ns,
x"00000000" AFTER 14740 ns,
x"EE6B276F" AFTER 14760 ns,
x"00000000" AFTER 14780 ns,
x"EE6B276B" AFTER 14800 ns,
x"00000000" AFTER 14820 ns,
x"EE6B2767" AFTER 14840 ns,
x"00000000" AFTER 14860 ns,
x"EE6B2763" AFTER 14880 ns,
x"00000000" AFTER 14900 ns,
x"EE6B275F" AFTER 14920 ns,
x"00000000" AFTER 14940 ns,
x"EE6B275B" AFTER 14960 ns,
x"00000000" AFTER 14980 ns,
x"EE6B2757" AFTER 15000 ns,
x"00000000" AFTER 15020 ns,
x"EE6B2753" AFTER 15040 ns,
x"00000000" AFTER 15060 ns,
x"EE6B274F" AFTER 15080 ns,
x"00000000" AFTER 15100 ns,
x"EE6B274B" AFTER 15120 ns,
x"00000000" AFTER 15140 ns,
x"EE6B2747" AFTER 15160 ns,
x"00000000" AFTER 15180 ns,
x"EE6B2743" AFTER 15200 ns,
x"00000000" AFTER 15220 ns,
x"EE6B273F" AFTER 15240 ns,
x"00000000" AFTER 15260 ns,
x"EE6B273B" AFTER 15280 ns,
x"00000000" AFTER 15300 ns,
x"EE6B2737" AFTER 15320 ns,
x"00000000" AFTER 15340 ns,
x"EE6B2733" AFTER 15360 ns,
x"00000000" AFTER 15380 ns,
x"EE6B272F" AFTER 15400 ns,
x"00000000" AFTER 15420 ns,
x"EE6B272B" AFTER 15440 ns,
x"00000000" AFTER 15460 ns,
x"EE6B2727" AFTER 15480 ns,
x"00000000" AFTER 15500 ns,
x"EE6B2723" AFTER 15520 ns,
x"00000000" AFTER 15540 ns,
x"EE6B271F" AFTER 15560 ns,
x"00000000" AFTER 15580 ns,
x"EE6B271B" AFTER 15600 ns,
x"00000000" AFTER 15620 ns,
x"EE6B2717" AFTER 15640 ns,
x"00000000" AFTER 15660 ns,
x"EE6B2713" AFTER 15680 ns,
x"00000000" AFTER 15700 ns,
x"EE6B270F" AFTER 15720 ns,
x"00000000" AFTER 15740 ns,
x"EE6B270B" AFTER 15760 ns,
x"00000000" AFTER 15780 ns,
x"EE6B2707" AFTER 15800 ns,
x"00000000" AFTER 15820 ns,
x"EE6B2703" AFTER 15840 ns,
x"00000000" AFTER 15860 ns,
x"EE6B26FF" AFTER 15880 ns,
x"00000000" AFTER 15900 ns,
x"EE6B26FB" AFTER 15920 ns,
x"00000000" AFTER 15940 ns,
x"EE6B26F7" AFTER 15960 ns,
x"00000000" AFTER 15980 ns,
x"EE6B26F3" AFTER 16000 ns,
x"00000000" AFTER 16020 ns,
x"EE6B26EF" AFTER 16040 ns,
x"00000000" AFTER 16060 ns,
x"EE6B26EB" AFTER 16080 ns,
x"00000000" AFTER 16100 ns,
x"EE6B26E7" AFTER 16120 ns,
x"00000000" AFTER 16140 ns,
x"EE6B26E3" AFTER 16160 ns,
x"00000000" AFTER 16180 ns,
x"EE6B26DF" AFTER 16200 ns,
x"00000000" AFTER 16220 ns,
x"EE6B26DB" AFTER 16240 ns,
x"00000000" AFTER 16260 ns,
x"EE6B26D7" AFTER 16280 ns,
x"00000000" AFTER 16300 ns,
x"EE6B26D3" AFTER 16320 ns,
x"00000000" AFTER 16340 ns,
x"EE6B26CF" AFTER 16360 ns,
x"00000000" AFTER 16380 ns,
x"EE6B26CB" AFTER 16400 ns,
x"00000000" AFTER 16420 ns,
x"EE6B26C7" AFTER 16440 ns,
x"00000000" AFTER 16460 ns,
x"EE6B26C3" AFTER 16480 ns,
x"00000000" AFTER 16500 ns,
x"EE6B26BF" AFTER 16520 ns,
x"00000000" AFTER 16540 ns,
x"EE6B26BB" AFTER 16560 ns,
x"00000000" AFTER 16580 ns,
x"EE6B26B7" AFTER 16600 ns,
x"00000000" AFTER 16620 ns,
x"EE6B26B3" AFTER 16640 ns,
x"00000000" AFTER 16660 ns,
x"EE6B26AF" AFTER 16680 ns,
x"00000000" AFTER 16700 ns,
x"EE6B26AB" AFTER 16720 ns,
x"00000000" AFTER 16740 ns,
x"EE6B26A7" AFTER 16760 ns,
x"00000000" AFTER 16780 ns,
x"EE6B26A3" AFTER 16800 ns,
x"00000000" AFTER 16820 ns,
x"EE6B269F" AFTER 16840 ns,
x"00000000" AFTER 16860 ns,
x"EE6B269B" AFTER 16880 ns,
x"00000000" AFTER 16900 ns,
x"EE6B2697" AFTER 16920 ns,
x"00000000" AFTER 16940 ns,
x"EE6B2693" AFTER 16960 ns,
x"00000000" AFTER 16980 ns,
x"EE6B268F" AFTER 17000 ns,
x"00000000" AFTER 17020 ns,
x"EE6B268B" AFTER 17040 ns,
x"00000000" AFTER 17060 ns,
x"EE6B2687" AFTER 17080 ns,
x"00000000" AFTER 17100 ns,
x"EE6B2683" AFTER 17120 ns,
x"00000000" AFTER 17140 ns,
x"EE6B267F" AFTER 17160 ns,
x"00000000" AFTER 17180 ns,
x"EE6B267B" AFTER 17200 ns,
x"00000000" AFTER 17220 ns,
x"EE6B2677" AFTER 17240 ns,
x"00000000" AFTER 17260 ns,
x"EE6B2673" AFTER 17280 ns,
x"00000000" AFTER 17300 ns,
x"EE6B266F" AFTER 17320 ns,
x"00000000" AFTER 17340 ns,
x"EE6B266B" AFTER 17360 ns,
x"00000000" AFTER 17380 ns,
x"EE6B2667" AFTER 17400 ns,
x"00000000" AFTER 17420 ns,
x"EE6B2663" AFTER 17440 ns,
x"00000000" AFTER 17460 ns,
x"EE6B265F" AFTER 17480 ns,
x"00000000" AFTER 17500 ns,
x"EE6B265B" AFTER 17520 ns,
x"00000000" AFTER 17540 ns,
x"EE6B2657" AFTER 17560 ns,
x"00000000" AFTER 17580 ns,
x"EE6B2653" AFTER 17600 ns,
x"00000000" AFTER 17620 ns,
x"EE6B264F" AFTER 17640 ns,
x"00000000" AFTER 17660 ns,
x"EE6B264B" AFTER 17680 ns,
x"00000000" AFTER 17700 ns,
x"EE6B2647" AFTER 17720 ns,
x"00000000" AFTER 17740 ns,
x"EE6B2643" AFTER 17760 ns,
x"00000000" AFTER 17780 ns,
x"EE6B263F" AFTER 17800 ns,
x"00000000" AFTER 17820 ns,
x"EE6B263B" AFTER 17840 ns,
x"00000000" AFTER 17860 ns,
x"EE6B2637" AFTER 17880 ns,
x"00000000" AFTER 17900 ns,
x"EE6B2633" AFTER 17920 ns,
x"00000000" AFTER 17940 ns,
x"EE6B262F" AFTER 17960 ns,
x"00000000" AFTER 17980 ns,
x"EE6B262B" AFTER 18000 ns,
x"00000000" AFTER 18020 ns,
x"EE6B2627" AFTER 18040 ns,
x"00000000" AFTER 18060 ns,
x"EE6B2623" AFTER 18080 ns,
x"00000000" AFTER 18100 ns,
x"EE6B261F" AFTER 18120 ns,
x"00000000" AFTER 18140 ns,
x"EE6B261B" AFTER 18160 ns,
x"00000000" AFTER 18180 ns,
x"EE6B2617" AFTER 18200 ns,
x"00000000" AFTER 18220 ns,
x"EE6B2613" AFTER 18240 ns,
x"00000000" AFTER 18260 ns,
x"EE6B260F" AFTER 18280 ns,
x"00000000" AFTER 18300 ns,
x"EE6B260B" AFTER 18320 ns,
x"00000000" AFTER 18340 ns,
x"EE6B2607" AFTER 18360 ns,
x"00000000" AFTER 18380 ns,
x"EE6B2603" AFTER 18400 ns,
x"00000000" AFTER 18420 ns,
x"EE6B25FF" AFTER 18440 ns,
x"00000000" AFTER 18460 ns,
x"EE6B25FB" AFTER 18480 ns,
x"00000000" AFTER 18500 ns,
x"EE6B25F7" AFTER 18520 ns,
x"00000000" AFTER 18540 ns,
x"EE6B25F3" AFTER 18560 ns,
x"00000000" AFTER 18580 ns,
x"EE6B25EF" AFTER 18600 ns,
x"00000000" AFTER 18620 ns,
x"EE6B25EB" AFTER 18640 ns,
x"00000000" AFTER 18660 ns,
x"EE6B25E7" AFTER 18680 ns,
x"00000000" AFTER 18700 ns,
x"EE6B25E3" AFTER 18720 ns,
x"00000000" AFTER 18740 ns,
x"EE6B25DF" AFTER 18760 ns,
x"00000000" AFTER 18780 ns,
x"EE6B25DB" AFTER 18800 ns,
x"00000000" AFTER 18820 ns,
x"EE6B25D7" AFTER 18840 ns,
x"00000000" AFTER 18860 ns,
x"EE6B25D3" AFTER 18880 ns,
x"00000000" AFTER 18900 ns,
x"EE6B25CF" AFTER 18920 ns,
x"00000000" AFTER 18940 ns,
x"EE6B25CB" AFTER 18960 ns,
x"00000000" AFTER 18980 ns,
x"EE6B25C7" AFTER 19000 ns,
x"00000000" AFTER 19020 ns,
x"EE6B25C3" AFTER 19040 ns,
x"00000000" AFTER 19060 ns,
x"EE6B25BF" AFTER 19080 ns,
x"00000000" AFTER 19100 ns,
x"EE6B25BB" AFTER 19120 ns,
x"00000000" AFTER 19140 ns,
x"EE6B25B7" AFTER 19160 ns,
x"00000000" AFTER 19180 ns,
x"EE6B25B3" AFTER 19200 ns,
x"00000000" AFTER 19220 ns,
x"EE6B25AF" AFTER 19240 ns,
x"00000000" AFTER 19260 ns,
x"EE6B25AB" AFTER 19280 ns,
x"00000000" AFTER 19300 ns,
x"EE6B25A7" AFTER 19320 ns,
x"00000000" AFTER 19340 ns,
x"EE6B25A3" AFTER 19360 ns,
x"00000000" AFTER 19380 ns,
x"EE6B259F" AFTER 19400 ns,
x"00000000" AFTER 19420 ns,
x"EE6B259B" AFTER 19440 ns,
x"00000000" AFTER 19460 ns,
x"EE6B2597" AFTER 19480 ns,
x"00000000" AFTER 19500 ns,
x"EE6B2593" AFTER 19520 ns,
x"00000000" AFTER 19540 ns,
x"EE6B258F" AFTER 19560 ns,
x"00000000" AFTER 19580 ns,
x"EE6B258B" AFTER 19600 ns,
x"00000000" AFTER 19620 ns,
x"EE6B2587" AFTER 19640 ns,
x"00000000" AFTER 19660 ns,
x"EE6B2583" AFTER 19680 ns,
x"00000000" AFTER 19700 ns,
x"EE6B257F" AFTER 19720 ns,
x"00000000" AFTER 19740 ns,
x"EE6B257B" AFTER 19760 ns,
x"00000000" AFTER 19780 ns,
x"EE6B2577" AFTER 19800 ns,
x"00000000" AFTER 19820 ns,
x"EE6B2573" AFTER 19840 ns,
x"00000000" AFTER 19860 ns,
x"EE6B256F" AFTER 19880 ns,
x"00000000" AFTER 19900 ns,
x"EE6B256B" AFTER 19920 ns,
x"00000000" AFTER 19940 ns,
x"EE6B256F" AFTER 19960 ns,
x"00000000" AFTER 19980 ns,
x"EE6B2573" AFTER 20000 ns,
x"00000000" AFTER 20020 ns,
x"EE6B2577" AFTER 20040 ns,
x"00000000" AFTER 20060 ns,
x"EE6B257B" AFTER 20080 ns,
x"00000000" AFTER 20100 ns,
x"EE6B257F" AFTER 20120 ns,
x"00000000" AFTER 20140 ns,
x"EE6B2583" AFTER 20160 ns,
x"00000000" AFTER 20180 ns,
x"EE6B2587" AFTER 20200 ns,
x"00000000" AFTER 20220 ns,
x"EE6B258B" AFTER 20240 ns,
x"00000000" AFTER 20260 ns,
x"EE6B258F" AFTER 20280 ns,
x"00000000" AFTER 20300 ns,
x"EE6B2593" AFTER 20320 ns,
x"00000000" AFTER 20340 ns,
x"EE6B2597" AFTER 20360 ns,
x"00000000" AFTER 20380 ns,
x"EE6B259B" AFTER 20400 ns,
x"00000000" AFTER 20420 ns,
x"EE6B259F" AFTER 20440 ns,
x"00000000" AFTER 20460 ns,
x"EE6B25A3" AFTER 20480 ns,
x"00000000" AFTER 20500 ns,
x"EE6B25A7" AFTER 20520 ns,
x"00000000" AFTER 20540 ns,
x"EE6B25AB" AFTER 20560 ns,
x"00000000" AFTER 20580 ns,
x"EE6B25AF" AFTER 20600 ns,
x"00000000" AFTER 20620 ns,
x"EE6B25B3" AFTER 20640 ns,
x"00000000" AFTER 20660 ns,
x"EE6B25B7" AFTER 20680 ns,
x"00000000" AFTER 20700 ns,
x"EE6B25BB" AFTER 20720 ns,
x"00000000" AFTER 20740 ns,
x"EE6B25BF" AFTER 20760 ns,
x"00000000" AFTER 20780 ns,
x"EE6B25C3" AFTER 20800 ns,
x"00000000" AFTER 20820 ns,
x"EE6B25C7" AFTER 20840 ns,
x"00000000" AFTER 20860 ns,
x"EE6B25CB" AFTER 20880 ns,
x"00000000" AFTER 20900 ns,
x"EE6B25CF" AFTER 20920 ns,
x"00000000" AFTER 20940 ns,
x"EE6B25D3" AFTER 20960 ns,
x"00000000" AFTER 20980 ns,
x"EE6B25D7" AFTER 21000 ns,
x"00000000" AFTER 21020 ns,
x"EE6B25DB" AFTER 21040 ns,
x"00000000" AFTER 21060 ns,
x"EE6B25DF" AFTER 21080 ns,
x"00000000" AFTER 21100 ns,
x"EE6B25E3" AFTER 21120 ns,
x"00000000" AFTER 21140 ns,
x"EE6B25E7" AFTER 21160 ns,
x"00000000" AFTER 21180 ns,
x"EE6B25EB" AFTER 21200 ns,
x"00000000" AFTER 21220 ns,
x"EE6B25EF" AFTER 21240 ns,
x"00000000" AFTER 21260 ns,
x"EE6B25F3" AFTER 21280 ns,
x"00000000" AFTER 21300 ns,
x"EE6B25F7" AFTER 21320 ns,
x"00000000" AFTER 21340 ns,
x"EE6B25FB" AFTER 21360 ns,
x"00000000" AFTER 21380 ns,
x"EE6B25FF" AFTER 21400 ns,
x"00000000" AFTER 21420 ns,
x"EE6B2603" AFTER 21440 ns,
x"00000000" AFTER 21460 ns,
x"EE6B2607" AFTER 21480 ns,
x"00000000" AFTER 21500 ns,
x"EE6B260B" AFTER 21520 ns,
x"00000000" AFTER 21540 ns,
x"EE6B260F" AFTER 21560 ns,
x"00000000" AFTER 21580 ns,
x"EE6B2613" AFTER 21600 ns,
x"00000000" AFTER 21620 ns,
x"EE6B2617" AFTER 21640 ns,
x"00000000" AFTER 21660 ns,
x"EE6B261B" AFTER 21680 ns,
x"00000000" AFTER 21700 ns,
x"EE6B261F" AFTER 21720 ns,
x"00000000" AFTER 21740 ns,
x"EE6B2623" AFTER 21760 ns,
x"00000000" AFTER 21780 ns,
x"EE6B2627" AFTER 21800 ns,
x"00000000" AFTER 21820 ns,
x"EE6B262B" AFTER 21840 ns,
x"00000000" AFTER 21860 ns,
x"EE6B262F" AFTER 21880 ns,
x"00000000" AFTER 21900 ns,
x"EE6B2633" AFTER 21920 ns,
x"00000000" AFTER 21940 ns,
x"EE6B2637" AFTER 21960 ns,
x"00000000" AFTER 21980 ns,
x"EE6B263B" AFTER 22000 ns,
x"00000000" AFTER 22020 ns,
x"EE6B263F" AFTER 22040 ns,
x"00000000" AFTER 22060 ns,
x"EE6B2643" AFTER 22080 ns,
x"00000000" AFTER 22100 ns,
x"EE6B2647" AFTER 22120 ns,
x"00000000" AFTER 22140 ns,
x"EE6B264B" AFTER 22160 ns,
x"00000000" AFTER 22180 ns,
x"EE6B264F" AFTER 22200 ns,
x"00000000" AFTER 22220 ns,
x"EE6B2653" AFTER 22240 ns,
x"00000000" AFTER 22260 ns,
x"EE6B2657" AFTER 22280 ns,
x"00000000" AFTER 22300 ns,
x"EE6B265B" AFTER 22320 ns,
x"00000000" AFTER 22340 ns,
x"EE6B265F" AFTER 22360 ns,
x"00000000" AFTER 22380 ns,
x"EE6B2663" AFTER 22400 ns,
x"00000000" AFTER 22420 ns,
x"EE6B2667" AFTER 22440 ns,
x"00000000" AFTER 22460 ns,
x"EE6B266B" AFTER 22480 ns,
x"00000000" AFTER 22500 ns,
x"EE6B266F" AFTER 22520 ns,
x"00000000" AFTER 22540 ns,
x"EE6B2673" AFTER 22560 ns,
x"00000000" AFTER 22580 ns,
x"EE6B2677" AFTER 22600 ns,
x"00000000" AFTER 22620 ns,
x"EE6B267B" AFTER 22640 ns,
x"00000000" AFTER 22660 ns,
x"EE6B267F" AFTER 22680 ns,
x"00000000" AFTER 22700 ns,
x"EE6B2683" AFTER 22720 ns,
x"00000000" AFTER 22740 ns,
x"EE6B2687" AFTER 22760 ns,
x"00000000" AFTER 22780 ns,
x"EE6B268B" AFTER 22800 ns,
x"00000000" AFTER 22820 ns,
x"EE6B268F" AFTER 22840 ns,
x"00000000" AFTER 22860 ns,
x"EE6B2693" AFTER 22880 ns,
x"00000000" AFTER 22900 ns,
x"EE6B2697" AFTER 22920 ns,
x"00000000" AFTER 22940 ns,
x"EE6B269B" AFTER 22960 ns,
x"00000000" AFTER 22980 ns,
x"EE6B269F" AFTER 23000 ns,
x"00000000" AFTER 23020 ns,
x"EE6B26A3" AFTER 23040 ns,
x"00000000" AFTER 23060 ns,
x"EE6B26A7" AFTER 23080 ns,
x"00000000" AFTER 23100 ns,
x"EE6B26AB" AFTER 23120 ns,
x"00000000" AFTER 23140 ns,
x"EE6B26AF" AFTER 23160 ns,
x"00000000" AFTER 23180 ns,
x"EE6B26B3" AFTER 23200 ns,
x"00000000" AFTER 23220 ns,
x"EE6B26B7" AFTER 23240 ns,
x"00000000" AFTER 23260 ns,
x"EE6B26BB" AFTER 23280 ns,
x"00000000" AFTER 23300 ns,
x"EE6B26BF" AFTER 23320 ns,
x"00000000" AFTER 23340 ns,
x"EE6B26C3" AFTER 23360 ns,
x"00000000" AFTER 23380 ns,
x"EE6B26C7" AFTER 23400 ns,
x"00000000" AFTER 23420 ns,
x"EE6B26CB" AFTER 23440 ns,
x"00000000" AFTER 23460 ns,
x"EE6B26CF" AFTER 23480 ns,
x"00000000" AFTER 23500 ns,
x"EE6B26D3" AFTER 23520 ns,
x"00000000" AFTER 23540 ns,
x"EE6B26D7" AFTER 23560 ns,
x"00000000" AFTER 23580 ns,
x"EE6B26DB" AFTER 23600 ns,
x"00000000" AFTER 23620 ns,
x"EE6B26DF" AFTER 23640 ns,
x"00000000" AFTER 23660 ns,
x"EE6B26E3" AFTER 23680 ns,
x"00000000" AFTER 23700 ns,
x"EE6B26E7" AFTER 23720 ns,
x"00000000" AFTER 23740 ns,
x"EE6B26EB" AFTER 23760 ns,
x"00000000" AFTER 23780 ns,
x"EE6B26EF" AFTER 23800 ns,
x"00000000" AFTER 23820 ns,
x"EE6B26F3" AFTER 23840 ns,
x"00000000" AFTER 23860 ns,
x"EE6B26F7" AFTER 23880 ns,
x"00000000" AFTER 23900 ns,
x"EE6B26FB" AFTER 23920 ns,
x"00000000" AFTER 23940 ns,
x"EE6B26FF" AFTER 23960 ns,
x"00000000" AFTER 23980 ns,
x"EE6B2703" AFTER 24000 ns,
x"00000000" AFTER 24020 ns,
x"EE6B2707" AFTER 24040 ns,
x"00000000" AFTER 24060 ns,
x"EE6B270B" AFTER 24080 ns,
x"00000000" AFTER 24100 ns,
x"EE6B270F" AFTER 24120 ns,
x"00000000" AFTER 24140 ns,
x"EE6B2713" AFTER 24160 ns,
x"00000000" AFTER 24180 ns,
x"EE6B2717" AFTER 24200 ns,
x"00000000" AFTER 24220 ns,
x"EE6B271B" AFTER 24240 ns,
x"00000000" AFTER 24260 ns,
x"EE6B271F" AFTER 24280 ns,
x"00000000" AFTER 24300 ns,
x"EE6B2723" AFTER 24320 ns,
x"00000000" AFTER 24340 ns,
x"EE6B2727" AFTER 24360 ns,
x"00000000" AFTER 24380 ns,
x"EE6B272B" AFTER 24400 ns,
x"00000000" AFTER 24420 ns,
x"EE6B272F" AFTER 24440 ns,
x"00000000" AFTER 24460 ns,
x"EE6B2733" AFTER 24480 ns,
x"00000000" AFTER 24500 ns,
x"EE6B2737" AFTER 24520 ns,
x"00000000" AFTER 24540 ns,
x"EE6B273B" AFTER 24560 ns,
x"00000000" AFTER 24580 ns,
x"EE6B273F" AFTER 24600 ns,
x"00000000" AFTER 24620 ns,
x"EE6B2743" AFTER 24640 ns,
x"00000000" AFTER 24660 ns,
x"EE6B2747" AFTER 24680 ns,
x"00000000" AFTER 24700 ns,
x"EE6B274B" AFTER 24720 ns,
x"00000000" AFTER 24740 ns,
x"EE6B274F" AFTER 24760 ns,
x"00000000" AFTER 24780 ns,
x"EE6B2753" AFTER 24800 ns,
x"00000000" AFTER 24820 ns,
x"EE6B2757" AFTER 24840 ns,
x"00000000" AFTER 24860 ns,
x"EE6B275B" AFTER 24880 ns,
x"00000000" AFTER 24900 ns,
x"EE6B275F" AFTER 24920 ns,
x"00000000" AFTER 24940 ns,
x"EE6B2763" AFTER 24960 ns,
x"00000000" AFTER 24980 ns,
x"EE6B2767" AFTER 25000 ns,
x"00000000" AFTER 25020 ns,
x"EE6B276B" AFTER 25040 ns,
x"00000000" AFTER 25060 ns,
x"EE6B276F" AFTER 25080 ns,
x"00000000" AFTER 25100 ns,
x"EE6B2773" AFTER 25120 ns,
x"00000000" AFTER 25140 ns,
x"EE6B2777" AFTER 25160 ns,
x"00000000" AFTER 25180 ns,
x"EE6B277B" AFTER 25200 ns,
x"00000000" AFTER 25220 ns,
x"EE6B277F" AFTER 25240 ns,
x"00000000" AFTER 25260 ns,
x"EE6B2783" AFTER 25280 ns,
x"00000000" AFTER 25300 ns,
x"EE6B2787" AFTER 25320 ns,
x"00000000" AFTER 25340 ns,
x"EE6B278B" AFTER 25360 ns,
x"00000000" AFTER 25380 ns,
x"EE6B278F" AFTER 25400 ns,
x"00000000" AFTER 25420 ns,
x"EE6B2793" AFTER 25440 ns,
x"00000000" AFTER 25460 ns,
x"EE6B2797" AFTER 25480 ns,
x"00000000" AFTER 25500 ns,
x"EE6B279B" AFTER 25520 ns,
x"00000000" AFTER 25540 ns,
x"EE6B279F" AFTER 25560 ns,
x"00000000" AFTER 25580 ns,
x"EE6B27A3" AFTER 25600 ns,
x"00000000" AFTER 25620 ns,
x"EE6B27A7" AFTER 25640 ns,
x"00000000" AFTER 25660 ns,
x"EE6B27AB" AFTER 25680 ns,
x"00000000" AFTER 25700 ns,
x"EE6B27AF" AFTER 25720 ns,
x"00000000" AFTER 25740 ns,
x"EE6B27B3" AFTER 25760 ns,
x"00000000" AFTER 25780 ns,
x"EE6B27B7" AFTER 25800 ns,
x"00000000" AFTER 25820 ns,
x"EE6B27BB" AFTER 25840 ns,
x"00000000" AFTER 25860 ns,
x"EE6B27BF" AFTER 25880 ns,
x"00000000" AFTER 25900 ns,
x"EE6B27C3" AFTER 25920 ns,
x"00000000" AFTER 25940 ns,
x"EE6B27C7" AFTER 25960 ns,
x"00000000" AFTER 25980 ns,
x"EE6B27CB" AFTER 26000 ns,
x"00000000" AFTER 26020 ns,
x"EE6B27CF" AFTER 26040 ns,
x"00000000" AFTER 26060 ns,
x"EE6B27D3" AFTER 26080 ns,
x"00000000" AFTER 26100 ns,
x"EE6B27D7" AFTER 26120 ns,
x"00000000" AFTER 26140 ns,
x"EE6B27DB" AFTER 26160 ns,
x"00000000" AFTER 26180 ns,
x"EE6B27DF" AFTER 26200 ns,
x"00000000" AFTER 26220 ns,
x"EE6B27E3" AFTER 26240 ns,
x"00000000" AFTER 26260 ns,
x"EE6B27E7" AFTER 26280 ns,
x"00000000" AFTER 26300 ns,
x"EE6B27EB" AFTER 26320 ns,
x"00000000" AFTER 26340 ns,
x"EE6B27EF" AFTER 26360 ns,
x"00000000" AFTER 26380 ns,
x"EE6B27F3" AFTER 26400 ns,
x"00000000" AFTER 26420 ns,
x"EE6B27F7" AFTER 26440 ns,
x"00000000" AFTER 26460 ns,
x"EE6B27FB" AFTER 26480 ns,
x"00000000" AFTER 26500 ns,
x"EE6B27FF" AFTER 26520 ns,
x"00000000" AFTER 26540 ns,
x"EE6B2803" AFTER 26560 ns,
x"00000000" AFTER 26580 ns,
x"EE6B2807" AFTER 26600 ns,
x"00000000" AFTER 26620 ns,
x"EE6B280B" AFTER 26640 ns,
x"00000000" AFTER 26660 ns,
x"EE6B280F" AFTER 26680 ns,
x"00000000" AFTER 26700 ns,
x"EE6B2813" AFTER 26720 ns,
x"00000000" AFTER 26740 ns,
x"EE6B2817" AFTER 26760 ns,
x"00000000" AFTER 26780 ns,
x"EE6B281B" AFTER 26800 ns,
x"00000000" AFTER 26820 ns,
x"EE6B281F" AFTER 26840 ns,
x"00000000" AFTER 26860 ns,
x"EE6B2823" AFTER 26880 ns,
x"00000000" AFTER 26900 ns,
x"EE6B2827" AFTER 26920 ns,
x"00000000" AFTER 26940 ns,
x"EE6B282B" AFTER 26960 ns,
x"00000000" AFTER 26980 ns,
x"EE6B282F" AFTER 27000 ns,
x"00000000" AFTER 27020 ns,
x"EE6B2833" AFTER 27040 ns,
x"00000000" AFTER 27060 ns,
x"EE6B2837" AFTER 27080 ns,
x"00000000" AFTER 27100 ns,
x"EE6B283B" AFTER 27120 ns,
x"00000000" AFTER 27140 ns,
x"EE6B283F" AFTER 27160 ns,
x"00000000" AFTER 27180 ns,
x"EE6B2843" AFTER 27200 ns,
x"00000000" AFTER 27220 ns,
x"EE6B2847" AFTER 27240 ns,
x"00000000" AFTER 27260 ns,
x"EE6B284B" AFTER 27280 ns,
x"00000000" AFTER 27300 ns,
x"EE6B284F" AFTER 27320 ns,
x"00000000" AFTER 27340 ns,
x"EE6B2853" AFTER 27360 ns,
x"00000000" AFTER 27380 ns,
x"EE6B2857" AFTER 27400 ns,
x"00000000" AFTER 27420 ns,
x"EE6B285B" AFTER 27440 ns,
x"00000000" AFTER 27460 ns,
x"EE6B285F" AFTER 27480 ns,
x"00000000" AFTER 27500 ns,
x"EE6B2863" AFTER 27520 ns,
x"00000000" AFTER 27540 ns,
x"EE6B2867" AFTER 27560 ns,
x"00000000" AFTER 27580 ns,
x"EE6B286B" AFTER 27600 ns,
x"00000000" AFTER 27620 ns,
x"EE6B286F" AFTER 27640 ns,
x"00000000" AFTER 27660 ns,
x"EE6B2873" AFTER 27680 ns,
x"00000000" AFTER 27700 ns,
x"EE6B2877" AFTER 27720 ns,
x"00000000" AFTER 27740 ns,
x"EE6B287B" AFTER 27760 ns,
x"00000000" AFTER 27780 ns,
x"EE6B287F" AFTER 27800 ns,
x"00000000" AFTER 27820 ns,
x"EE6B2883" AFTER 27840 ns,
x"00000000" AFTER 27860 ns,
x"EE6B2887" AFTER 27880 ns,
x"00000000" AFTER 27900 ns,
x"EE6B288B" AFTER 27920 ns,
x"00000000" AFTER 27940 ns,
x"EE6B288F" AFTER 27960 ns,
x"00000000" AFTER 27980 ns,
x"EE6B2893" AFTER 28000 ns,
x"00000000" AFTER 28020 ns,
x"EE6B2897" AFTER 28040 ns,
x"00000000" AFTER 28060 ns,
x"EE6B289B" AFTER 28080 ns,
x"00000000" AFTER 28100 ns,
x"EE6B289F" AFTER 28120 ns,
x"00000000" AFTER 28140 ns,
x"EE6B28A3" AFTER 28160 ns,
x"00000000" AFTER 28180 ns,
x"EE6B28A7" AFTER 28200 ns,
x"00000000" AFTER 28220 ns,
x"EE6B28AB" AFTER 28240 ns,
x"00000000" AFTER 28260 ns,
x"EE6B28AF" AFTER 28280 ns,
x"00000000" AFTER 28300 ns,
x"EE6B28B3" AFTER 28320 ns,
x"00000000" AFTER 28340 ns,
x"EE6B28B7" AFTER 28360 ns,
x"00000000" AFTER 28380 ns,
x"EE6B28BB" AFTER 28400 ns,
x"00000000" AFTER 28420 ns,
x"EE6B28BF" AFTER 28440 ns,
x"00000000" AFTER 28460 ns,
x"EE6B28C3" AFTER 28480 ns,
x"00000000" AFTER 28500 ns,
x"EE6B28C7" AFTER 28520 ns,
x"00000000" AFTER 28540 ns,
x"EE6B28CB" AFTER 28560 ns,
x"00000000" AFTER 28580 ns,
x"EE6B28CF" AFTER 28600 ns,
x"00000000" AFTER 28620 ns,
x"EE6B28D3" AFTER 28640 ns,
x"00000000" AFTER 28660 ns,
x"EE6B28D7" AFTER 28680 ns,
x"00000000" AFTER 28700 ns,
x"EE6B28DB" AFTER 28720 ns,
x"00000000" AFTER 28740 ns,
x"EE6B28DF" AFTER 28760 ns,
x"00000000" AFTER 28780 ns,
x"EE6B28E3" AFTER 28800 ns,
x"00000000" AFTER 28820 ns,
x"EE6B28E7" AFTER 28840 ns,
x"00000000" AFTER 28860 ns,
x"EE6B28EB" AFTER 28880 ns,
x"00000000" AFTER 28900 ns,
x"EE6B28EF" AFTER 28920 ns,
x"00000000" AFTER 28940 ns,
x"EE6B28F3" AFTER 28960 ns,
x"00000000" AFTER 28980 ns,
x"EE6B28F7" AFTER 29000 ns,
x"00000000" AFTER 29020 ns,
x"EE6B28FB" AFTER 29040 ns,
x"00000000" AFTER 29060 ns,
x"EE6B28FF" AFTER 29080 ns,
x"00000000" AFTER 29100 ns,
x"EE6B2903" AFTER 29120 ns,
x"00000000" AFTER 29140 ns,
x"EE6B2907" AFTER 29160 ns,
x"00000000" AFTER 29180 ns,
x"EE6B290B" AFTER 29200 ns,
x"00000000" AFTER 29220 ns,
x"EE6B290F" AFTER 29240 ns,
x"00000000" AFTER 29260 ns,
x"EE6B2913" AFTER 29280 ns,
x"00000000" AFTER 29300 ns,
x"EE6B2917" AFTER 29320 ns,
x"00000000" AFTER 29340 ns,
x"EE6B291B" AFTER 29360 ns,
x"00000000" AFTER 29380 ns,
x"EE6B291F" AFTER 29400 ns,
x"00000000" AFTER 29420 ns,
x"EE6B2923" AFTER 29440 ns,
x"00000000" AFTER 29460 ns,
x"EE6B2927" AFTER 29480 ns,
x"00000000" AFTER 29500 ns,
x"EE6B292B" AFTER 29520 ns,
x"00000000" AFTER 29540 ns,
x"EE6B292F" AFTER 29560 ns,
x"00000000" AFTER 29580 ns,
x"EE6B2933" AFTER 29600 ns,
x"00000000" AFTER 29620 ns,
x"EE6B2937" AFTER 29640 ns,
x"00000000" AFTER 29660 ns,
x"EE6B293B" AFTER 29680 ns,
x"00000000" AFTER 29700 ns,
x"EE6B293F" AFTER 29720 ns,
x"00000000" AFTER 29740 ns,
x"EE6B2943" AFTER 29760 ns,
x"00000000" AFTER 29780 ns,
x"EE6B2947" AFTER 29800 ns,
x"00000000" AFTER 29820 ns,
x"EE6B294B" AFTER 29840 ns,
x"00000000" AFTER 29860 ns,
x"EE6B294F" AFTER 29880 ns,
x"00000000" AFTER 29900 ns,
x"EE6B2953" AFTER 29920 ns,
x"00000000" AFTER 29940 ns,
x"EE6B2957" AFTER 29960 ns,
x"00000000" AFTER 29980 ns,
x"EE6B295B" AFTER 30000 ns,
x"00000000" AFTER 30020 ns,
x"EE6B295F" AFTER 30040 ns,
x"00000000" AFTER 30060 ns,
x"EE6B2963" AFTER 30080 ns,
x"00000000" AFTER 30100 ns,
x"EE6B2967" AFTER 30120 ns,
x"00000000" AFTER 30140 ns,
x"EE6B296B" AFTER 30160 ns,
x"00000000" AFTER 30180 ns,
x"EE6B296F" AFTER 30200 ns,
x"00000000" AFTER 30220 ns,
x"EE6B2973" AFTER 30240 ns,
x"00000000" AFTER 30260 ns,
x"EE6B2977" AFTER 30280 ns,
x"00000000" AFTER 30300 ns,
x"EE6B297B" AFTER 30320 ns,
x"00000000" AFTER 30340 ns,
x"EE6B297F" AFTER 30360 ns,
x"00000000" AFTER 30380 ns,
x"EE6B2983" AFTER 30400 ns,
x"00000000" AFTER 30420 ns,
x"EE6B2987" AFTER 30440 ns,
x"00000000" AFTER 30460 ns,
x"EE6B298B" AFTER 30480 ns,
x"00000000" AFTER 30500 ns,
x"EE6B298F" AFTER 30520 ns,
x"00000000" AFTER 30540 ns,
x"EE6B2993" AFTER 30560 ns,
x"00000000" AFTER 30580 ns,
x"EE6B2997" AFTER 30600 ns,
x"00000000" AFTER 30620 ns,
x"EE6B299B" AFTER 30640 ns,
x"00000000" AFTER 30660 ns,
x"EE6B299F" AFTER 30680 ns,
x"00000000" AFTER 30700 ns,
x"EE6B29A3" AFTER 30720 ns,
x"00000000" AFTER 30740 ns,
x"EE6B29A7" AFTER 30760 ns,
x"00000000" AFTER 30780 ns,
x"EE6B29AB" AFTER 30800 ns,
x"00000000" AFTER 30820 ns,
x"EE6B29AF" AFTER 30840 ns,
x"00000000" AFTER 30860 ns,
x"EE6B29B3" AFTER 30880 ns,
x"00000000" AFTER 30900 ns,
x"EE6B29B7" AFTER 30920 ns,
x"00000000" AFTER 30940 ns,
x"EE6B29BB" AFTER 30960 ns;

MemoryOut <= x"00000000" AFTER 00020 ns,
x"00000534" AFTER 00040 ns,
x"00000000" AFTER 00060 ns,
x"00000530" AFTER 00080 ns,
x"00000000" AFTER 00100 ns,
x"0000052C" AFTER 00120 ns,
x"00000000" AFTER 00140 ns,
x"00000528" AFTER 00160 ns,
x"00000000" AFTER 00180 ns,
x"00000524" AFTER 00200 ns,
x"00000000" AFTER 00220 ns,
x"00000520" AFTER 00240 ns,
x"00000000" AFTER 00260 ns,
x"0000051C" AFTER 00280 ns,
x"00000000" AFTER 00300 ns,
x"00000518" AFTER 00320 ns,
x"00000000" AFTER 00340 ns,
x"00000514" AFTER 00360 ns,
x"00000000" AFTER 00380 ns,
x"00000510" AFTER 00400 ns,
x"00000000" AFTER 00420 ns,
x"0000050C" AFTER 00440 ns,
x"00000000" AFTER 00460 ns,
x"00000508" AFTER 00480 ns,
x"00000000" AFTER 00500 ns,
x"00000504" AFTER 00520 ns,
x"00000000" AFTER 00540 ns,
x"00000500" AFTER 00560 ns,
x"00000000" AFTER 00580 ns,
x"000004FC" AFTER 00600 ns,
x"00000000" AFTER 00620 ns,
x"000004F8" AFTER 00640 ns,
x"00000000" AFTER 00660 ns,
x"000004F4" AFTER 00680 ns,
x"00000000" AFTER 00700 ns,
x"000004F0" AFTER 00720 ns,
x"00000000" AFTER 00740 ns,
x"000004EC" AFTER 00760 ns,
x"00000000" AFTER 00780 ns,
x"000004E8" AFTER 00800 ns,
x"00000000" AFTER 00820 ns,
x"000004E4" AFTER 00840 ns,
x"00000000" AFTER 00860 ns,
x"000004E0" AFTER 00880 ns,
x"00000000" AFTER 00900 ns,
x"000004DC" AFTER 00920 ns,
x"00000000" AFTER 00940 ns,
x"000004D8" AFTER 00960 ns,
x"00000000" AFTER 00980 ns,
x"000004D4" AFTER 01000 ns,
x"00000000" AFTER 01020 ns,
x"000004D0" AFTER 01040 ns,
x"00000000" AFTER 01060 ns,
x"000004CC" AFTER 01080 ns,
x"00000000" AFTER 01100 ns,
x"000004C8" AFTER 01120 ns,
x"00000000" AFTER 01140 ns,
x"000004C4" AFTER 01160 ns,
x"00000000" AFTER 01180 ns,
x"000004C0" AFTER 01200 ns,
x"00000000" AFTER 01220 ns,
x"000004BC" AFTER 01240 ns,
x"00000000" AFTER 01260 ns,
x"000004B8" AFTER 01280 ns,
x"00000000" AFTER 01300 ns,
x"000004B4" AFTER 01320 ns,
x"00000000" AFTER 01340 ns,
x"000004B0" AFTER 01360 ns,
x"00000000" AFTER 01380 ns,
x"000004AC" AFTER 01400 ns,
x"00000000" AFTER 01420 ns,
x"000004A8" AFTER 01440 ns,
x"00000000" AFTER 01460 ns,
x"000004A4" AFTER 01480 ns,
x"00000000" AFTER 01500 ns,
x"000004A0" AFTER 01520 ns,
x"00000000" AFTER 01540 ns,
x"0000049C" AFTER 01560 ns,
x"00000000" AFTER 01580 ns,
x"00000498" AFTER 01600 ns,
x"00000000" AFTER 01620 ns,
x"00000494" AFTER 01640 ns,
x"00000000" AFTER 01660 ns,
x"00000490" AFTER 01680 ns,
x"00000000" AFTER 01700 ns,
x"0000048C" AFTER 01720 ns,
x"00000000" AFTER 01740 ns,
x"00000488" AFTER 01760 ns,
x"00000000" AFTER 01780 ns,
x"00000484" AFTER 01800 ns,
x"00000000" AFTER 01820 ns,
x"00000480" AFTER 01840 ns,
x"00000000" AFTER 01860 ns,
x"0000047C" AFTER 01880 ns,
x"00000000" AFTER 01900 ns,
x"00000478" AFTER 01920 ns,
x"00000000" AFTER 01940 ns,
x"00000474" AFTER 01960 ns,
x"00000000" AFTER 01980 ns,
x"00000470" AFTER 02000 ns,
x"00000000" AFTER 02020 ns,
x"0000046C" AFTER 02040 ns,
x"00000000" AFTER 02060 ns,
x"00000468" AFTER 02080 ns,
x"00000000" AFTER 02100 ns,
x"00000464" AFTER 02120 ns,
x"00000000" AFTER 02140 ns,
x"00000460" AFTER 02160 ns,
x"00000000" AFTER 02180 ns,
x"0000045C" AFTER 02200 ns,
x"00000000" AFTER 02220 ns,
x"00000458" AFTER 02240 ns,
x"00000000" AFTER 02260 ns,
x"00000454" AFTER 02280 ns,
x"00000000" AFTER 02300 ns,
x"00000450" AFTER 02320 ns,
x"00000000" AFTER 02340 ns,
x"0000044C" AFTER 02360 ns,
x"00000000" AFTER 02380 ns,
x"00000448" AFTER 02400 ns,
x"00000000" AFTER 02420 ns,
x"00000444" AFTER 02440 ns,
x"00000000" AFTER 02460 ns,
x"00000440" AFTER 02480 ns,
x"00000000" AFTER 02500 ns,
x"0000043C" AFTER 02520 ns,
x"00000000" AFTER 02540 ns,
x"00000438" AFTER 02560 ns,
x"00000000" AFTER 02580 ns,
x"00000434" AFTER 02600 ns,
x"00000000" AFTER 02620 ns,
x"00000430" AFTER 02640 ns,
x"00000000" AFTER 02660 ns,
x"0000042C" AFTER 02680 ns,
x"00000000" AFTER 02700 ns,
x"00000428" AFTER 02720 ns,
x"00000000" AFTER 02740 ns,
x"00000424" AFTER 02760 ns,
x"00000000" AFTER 02780 ns,
x"00000420" AFTER 02800 ns,
x"00000000" AFTER 02820 ns,
x"0000041C" AFTER 02840 ns,
x"00000000" AFTER 02860 ns,
x"00000418" AFTER 02880 ns,
x"00000000" AFTER 02900 ns,
x"00000414" AFTER 02920 ns,
x"00000000" AFTER 02940 ns,
x"00000410" AFTER 02960 ns,
x"00000000" AFTER 02980 ns,
x"0000040C" AFTER 03000 ns,
x"00000000" AFTER 03020 ns,
x"00000408" AFTER 03040 ns,
x"00000000" AFTER 03060 ns,
x"00000404" AFTER 03080 ns,
x"00000000" AFTER 03100 ns,
x"00000400" AFTER 03120 ns,
x"00000000" AFTER 03140 ns,
x"000003FC" AFTER 03160 ns,
x"00000000" AFTER 03180 ns,
x"000003F8" AFTER 03200 ns,
x"00000000" AFTER 03220 ns,
x"000003F4" AFTER 03240 ns,
x"00000000" AFTER 03260 ns,
x"000003F0" AFTER 03280 ns,
x"00000000" AFTER 03300 ns,
x"000003EC" AFTER 03320 ns,
x"00000000" AFTER 03340 ns,
x"000003E8" AFTER 03360 ns,
x"00000000" AFTER 03380 ns,
x"000003E4" AFTER 03400 ns,
x"00000000" AFTER 03420 ns,
x"000003E0" AFTER 03440 ns,
x"00000000" AFTER 03460 ns,
x"000003DC" AFTER 03480 ns,
x"00000000" AFTER 03500 ns,
x"000003D8" AFTER 03520 ns,
x"00000000" AFTER 03540 ns,
x"000003D4" AFTER 03560 ns,
x"00000000" AFTER 03580 ns,
x"000003D0" AFTER 03600 ns,
x"00000000" AFTER 03620 ns,
x"000003CC" AFTER 03640 ns,
x"00000000" AFTER 03660 ns,
x"000003C8" AFTER 03680 ns,
x"00000000" AFTER 03700 ns,
x"000003C4" AFTER 03720 ns,
x"00000000" AFTER 03740 ns,
x"000003C0" AFTER 03760 ns,
x"00000000" AFTER 03780 ns,
x"000003BC" AFTER 03800 ns,
x"00000000" AFTER 03820 ns,
x"000003B8" AFTER 03840 ns,
x"00000000" AFTER 03860 ns,
x"000003B4" AFTER 03880 ns,
x"00000000" AFTER 03900 ns,
x"000003B0" AFTER 03920 ns,
x"00000000" AFTER 03940 ns,
x"000003AC" AFTER 03960 ns,
x"00000000" AFTER 03980 ns,
x"000003A8" AFTER 04000 ns,
x"00000000" AFTER 04020 ns,
x"000003A4" AFTER 04040 ns,
x"00000000" AFTER 04060 ns,
x"000003A0" AFTER 04080 ns,
x"00000000" AFTER 04100 ns,
x"0000039C" AFTER 04120 ns,
x"00000000" AFTER 04140 ns,
x"00000398" AFTER 04160 ns,
x"00000000" AFTER 04180 ns,
x"00000394" AFTER 04200 ns,
x"00000000" AFTER 04220 ns,
x"00000390" AFTER 04240 ns,
x"00000000" AFTER 04260 ns,
x"0000038C" AFTER 04280 ns,
x"00000000" AFTER 04300 ns,
x"00000388" AFTER 04320 ns,
x"00000000" AFTER 04340 ns,
x"00000384" AFTER 04360 ns,
x"00000000" AFTER 04380 ns,
x"00000380" AFTER 04400 ns,
x"00000000" AFTER 04420 ns,
x"0000037C" AFTER 04440 ns,
x"00000000" AFTER 04460 ns,
x"00000378" AFTER 04480 ns,
x"00000000" AFTER 04500 ns,
x"00000374" AFTER 04520 ns,
x"00000000" AFTER 04540 ns,
x"00000370" AFTER 04560 ns,
x"00000000" AFTER 04580 ns,
x"0000036C" AFTER 04600 ns,
x"00000000" AFTER 04620 ns,
x"00000368" AFTER 04640 ns,
x"00000000" AFTER 04660 ns,
x"00000364" AFTER 04680 ns,
x"00000000" AFTER 04700 ns,
x"00000360" AFTER 04720 ns,
x"00000000" AFTER 04740 ns,
x"0000035C" AFTER 04760 ns,
x"00000000" AFTER 04780 ns,
x"00000358" AFTER 04800 ns,
x"00000000" AFTER 04820 ns,
x"00000354" AFTER 04840 ns,
x"00000000" AFTER 04860 ns,
x"00000350" AFTER 04880 ns,
x"00000000" AFTER 04900 ns,
x"0000034C" AFTER 04920 ns,
x"00000000" AFTER 04940 ns,
x"00000348" AFTER 04960 ns,
x"00000000" AFTER 04980 ns,
x"00000344" AFTER 05000 ns,
x"00000000" AFTER 05020 ns,
x"00000340" AFTER 05040 ns,
x"00000000" AFTER 05060 ns,
x"0000033C" AFTER 05080 ns,
x"00000000" AFTER 05100 ns,
x"00000338" AFTER 05120 ns,
x"00000000" AFTER 05140 ns,
x"00000334" AFTER 05160 ns,
x"00000000" AFTER 05180 ns,
x"00000330" AFTER 05200 ns,
x"00000000" AFTER 05220 ns,
x"0000032C" AFTER 05240 ns,
x"00000000" AFTER 05260 ns,
x"00000328" AFTER 05280 ns,
x"00000000" AFTER 05300 ns,
x"00000324" AFTER 05320 ns,
x"00000000" AFTER 05340 ns,
x"00000320" AFTER 05360 ns,
x"00000000" AFTER 05380 ns,
x"0000031C" AFTER 05400 ns,
x"00000000" AFTER 05420 ns,
x"00000318" AFTER 05440 ns,
x"00000000" AFTER 05460 ns,
x"00000314" AFTER 05480 ns,
x"00000000" AFTER 05500 ns,
x"00000310" AFTER 05520 ns,
x"00000000" AFTER 05540 ns,
x"0000030C" AFTER 05560 ns,
x"00000000" AFTER 05580 ns,
x"00000308" AFTER 05600 ns,
x"00000000" AFTER 05620 ns,
x"00000304" AFTER 05640 ns,
x"00000000" AFTER 05660 ns,
x"00000300" AFTER 05680 ns,
x"00000000" AFTER 05700 ns,
x"000002FC" AFTER 05720 ns,
x"00000000" AFTER 05740 ns,
x"000002F8" AFTER 05760 ns,
x"00000000" AFTER 05780 ns,
x"000002F4" AFTER 05800 ns,
x"00000000" AFTER 05820 ns,
x"000002F0" AFTER 05840 ns,
x"00000000" AFTER 05860 ns,
x"000002EC" AFTER 05880 ns,
x"00000000" AFTER 05900 ns,
x"000002E8" AFTER 05920 ns,
x"00000000" AFTER 05940 ns,
x"000002E4" AFTER 05960 ns,
x"00000000" AFTER 05980 ns,
x"000002E0" AFTER 06000 ns,
x"00000000" AFTER 06020 ns,
x"000002DC" AFTER 06040 ns,
x"00000000" AFTER 06060 ns,
x"000002D8" AFTER 06080 ns,
x"00000000" AFTER 06100 ns,
x"000002D4" AFTER 06120 ns,
x"00000000" AFTER 06140 ns,
x"000002D0" AFTER 06160 ns,
x"00000000" AFTER 06180 ns,
x"000002CC" AFTER 06200 ns,
x"00000000" AFTER 06220 ns,
x"000002C8" AFTER 06240 ns,
x"00000000" AFTER 06260 ns,
x"000002C4" AFTER 06280 ns,
x"00000000" AFTER 06300 ns,
x"000002C0" AFTER 06320 ns,
x"00000000" AFTER 06340 ns,
x"000002BC" AFTER 06360 ns,
x"00000000" AFTER 06380 ns,
x"000002B8" AFTER 06400 ns,
x"00000000" AFTER 06420 ns,
x"000002B4" AFTER 06440 ns,
x"00000000" AFTER 06460 ns,
x"000002B0" AFTER 06480 ns,
x"00000000" AFTER 06500 ns,
x"000002AC" AFTER 06520 ns,
x"00000000" AFTER 06540 ns,
x"000002A8" AFTER 06560 ns,
x"00000000" AFTER 06580 ns,
x"000002A4" AFTER 06600 ns,
x"00000000" AFTER 06620 ns,
x"000002A0" AFTER 06640 ns,
x"00000000" AFTER 06660 ns,
x"0000029C" AFTER 06680 ns,
x"00000000" AFTER 06700 ns,
x"00000298" AFTER 06720 ns,
x"00000000" AFTER 06740 ns,
x"00000294" AFTER 06760 ns,
x"00000000" AFTER 06780 ns,
x"00000290" AFTER 06800 ns,
x"00000000" AFTER 06820 ns,
x"0000028C" AFTER 06840 ns,
x"00000000" AFTER 06860 ns,
x"00000288" AFTER 06880 ns,
x"00000000" AFTER 06900 ns,
x"00000284" AFTER 06920 ns,
x"00000000" AFTER 06940 ns,
x"00000280" AFTER 06960 ns,
x"00000000" AFTER 06980 ns,
x"0000027C" AFTER 07000 ns,
x"00000000" AFTER 07020 ns,
x"00000278" AFTER 07040 ns,
x"00000000" AFTER 07060 ns,
x"00000274" AFTER 07080 ns,
x"00000000" AFTER 07100 ns,
x"00000270" AFTER 07120 ns,
x"00000000" AFTER 07140 ns,
x"0000026C" AFTER 07160 ns,
x"00000000" AFTER 07180 ns,
x"00000268" AFTER 07200 ns,
x"00000000" AFTER 07220 ns,
x"00000264" AFTER 07240 ns,
x"00000000" AFTER 07260 ns,
x"00000260" AFTER 07280 ns,
x"00000000" AFTER 07300 ns,
x"0000025C" AFTER 07320 ns,
x"00000000" AFTER 07340 ns,
x"00000258" AFTER 07360 ns,
x"00000000" AFTER 07380 ns,
x"00000254" AFTER 07400 ns,
x"00000000" AFTER 07420 ns,
x"00000250" AFTER 07440 ns,
x"00000000" AFTER 07460 ns,
x"0000024C" AFTER 07480 ns,
x"00000000" AFTER 07500 ns,
x"00000248" AFTER 07520 ns,
x"00000000" AFTER 07540 ns,
x"00000244" AFTER 07560 ns,
x"00000000" AFTER 07580 ns,
x"00000240" AFTER 07600 ns,
x"00000000" AFTER 07620 ns,
x"0000023C" AFTER 07640 ns,
x"00000000" AFTER 07660 ns,
x"00000238" AFTER 07680 ns,
x"00000000" AFTER 07700 ns,
x"00000234" AFTER 07720 ns,
x"00000000" AFTER 07740 ns,
x"00000230" AFTER 07760 ns,
x"00000000" AFTER 07780 ns,
x"0000022C" AFTER 07800 ns,
x"00000000" AFTER 07820 ns,
x"00000228" AFTER 07840 ns,
x"00000000" AFTER 07860 ns,
x"00000224" AFTER 07880 ns,
x"00000000" AFTER 07900 ns,
x"00000220" AFTER 07920 ns,
x"00000000" AFTER 07940 ns,
x"0000021C" AFTER 07960 ns,
x"00000000" AFTER 07980 ns,
x"00000218" AFTER 08000 ns,
x"00000000" AFTER 08020 ns,
x"00000214" AFTER 08040 ns,
x"00000000" AFTER 08060 ns,
x"00000210" AFTER 08080 ns,
x"00000000" AFTER 08100 ns,
x"0000020C" AFTER 08120 ns,
x"00000000" AFTER 08140 ns,
x"00000208" AFTER 08160 ns,
x"00000000" AFTER 08180 ns,
x"00000204" AFTER 08200 ns,
x"00000000" AFTER 08220 ns,
x"00000200" AFTER 08240 ns,
x"00000000" AFTER 08260 ns,
x"000001FC" AFTER 08280 ns,
x"00000000" AFTER 08300 ns,
x"000001F8" AFTER 08320 ns,
x"00000000" AFTER 08340 ns,
x"000001F4" AFTER 08360 ns,
x"00000000" AFTER 08380 ns,
x"000001F0" AFTER 08400 ns,
x"00000000" AFTER 08420 ns,
x"000001EC" AFTER 08440 ns,
x"00000000" AFTER 08460 ns,
x"000001E8" AFTER 08480 ns,
x"00000000" AFTER 08500 ns,
x"000001E4" AFTER 08520 ns,
x"00000000" AFTER 08540 ns,
x"000001E0" AFTER 08560 ns,
x"00000000" AFTER 08580 ns,
x"000001DC" AFTER 08600 ns,
x"00000000" AFTER 08620 ns,
x"000001D8" AFTER 08640 ns,
x"00000000" AFTER 08660 ns,
x"000001D4" AFTER 08680 ns,
x"00000000" AFTER 08700 ns,
x"000001D0" AFTER 08720 ns,
x"00000000" AFTER 08740 ns,
x"000001CC" AFTER 08760 ns,
x"00000000" AFTER 08780 ns,
x"000001C8" AFTER 08800 ns,
x"00000000" AFTER 08820 ns,
x"000001C4" AFTER 08840 ns,
x"00000000" AFTER 08860 ns,
x"000001C0" AFTER 08880 ns,
x"00000000" AFTER 08900 ns,
x"000001BC" AFTER 08920 ns,
x"00000000" AFTER 08940 ns,
x"000001B8" AFTER 08960 ns,
x"00000000" AFTER 08980 ns,
x"000001B4" AFTER 09000 ns,
x"00000000" AFTER 09020 ns,
x"000001B0" AFTER 09040 ns,
x"00000000" AFTER 09060 ns,
x"000001AC" AFTER 09080 ns,
x"00000000" AFTER 09100 ns,
x"000001A8" AFTER 09120 ns,
x"00000000" AFTER 09140 ns,
x"000001A4" AFTER 09160 ns,
x"00000000" AFTER 09180 ns,
x"000001A0" AFTER 09200 ns,
x"00000000" AFTER 09220 ns,
x"0000019C" AFTER 09240 ns,
x"00000000" AFTER 09260 ns,
x"00000198" AFTER 09280 ns,
x"00000000" AFTER 09300 ns,
x"00000194" AFTER 09320 ns,
x"00000000" AFTER 09340 ns,
x"00000190" AFTER 09360 ns,
x"00000000" AFTER 09380 ns,
x"0000018C" AFTER 09400 ns,
x"00000000" AFTER 09420 ns,
x"00000188" AFTER 09440 ns,
x"00000000" AFTER 09460 ns,
x"00000184" AFTER 09480 ns,
x"00000000" AFTER 09500 ns,
x"00000180" AFTER 09520 ns,
x"00000000" AFTER 09540 ns,
x"0000017C" AFTER 09560 ns,
x"00000000" AFTER 09580 ns,
x"00000178" AFTER 09600 ns,
x"00000000" AFTER 09620 ns,
x"00000174" AFTER 09640 ns,
x"00000000" AFTER 09660 ns,
x"00000170" AFTER 09680 ns,
x"00000000" AFTER 09700 ns,
x"0000016C" AFTER 09720 ns,
x"00000000" AFTER 09740 ns,
x"00000168" AFTER 09760 ns,
x"00000000" AFTER 09780 ns,
x"00000164" AFTER 09800 ns,
x"00000000" AFTER 09820 ns,
x"00000160" AFTER 09840 ns,
x"00000000" AFTER 09860 ns,
x"0000015C" AFTER 09880 ns,
x"00000000" AFTER 09900 ns,
x"00000158" AFTER 09920 ns,
x"00000000" AFTER 09940 ns,
x"00000154" AFTER 09960 ns,
x"00000000" AFTER 09980 ns,
x"00000150" AFTER 10000 ns,
x"00000000" AFTER 10020 ns,
x"0000014C" AFTER 10040 ns,
x"00000000" AFTER 10060 ns,
x"00000148" AFTER 10080 ns,
x"00000000" AFTER 10100 ns,
x"00000144" AFTER 10120 ns,
x"00000000" AFTER 10140 ns,
x"00000140" AFTER 10160 ns,
x"00000000" AFTER 10180 ns,
x"0000013C" AFTER 10200 ns,
x"00000000" AFTER 10220 ns,
x"00000138" AFTER 10240 ns,
x"00000000" AFTER 10260 ns,
x"00000134" AFTER 10280 ns,
x"00000000" AFTER 10300 ns,
x"00000130" AFTER 10320 ns,
x"00000000" AFTER 10340 ns,
x"0000012C" AFTER 10360 ns,
x"00000000" AFTER 10380 ns,
x"00000128" AFTER 10400 ns,
x"00000000" AFTER 10420 ns,
x"00000124" AFTER 10440 ns,
x"00000000" AFTER 10460 ns,
x"00000120" AFTER 10480 ns,
x"00000000" AFTER 10500 ns,
x"0000011C" AFTER 10520 ns,
x"00000000" AFTER 10540 ns,
x"00000118" AFTER 10560 ns,
x"00000000" AFTER 10580 ns,
x"00000114" AFTER 10600 ns,
x"00000000" AFTER 10620 ns,
x"00000110" AFTER 10640 ns,
x"00000000" AFTER 10660 ns,
x"0000010C" AFTER 10680 ns,
x"00000000" AFTER 10700 ns,
x"00000108" AFTER 10720 ns,
x"00000000" AFTER 10740 ns,
x"00000104" AFTER 10760 ns,
x"00000000" AFTER 10780 ns,
x"00000100" AFTER 10800 ns,
x"00000000" AFTER 10820 ns,
x"000000FC" AFTER 10840 ns,
x"00000000" AFTER 10860 ns,
x"000000F8" AFTER 10880 ns,
x"00000000" AFTER 10900 ns,
x"000000F4" AFTER 10920 ns,
x"00000000" AFTER 10940 ns,
x"000000F0" AFTER 10960 ns,
x"00000000" AFTER 10980 ns,
x"000000EC" AFTER 11000 ns,
x"00000000" AFTER 11020 ns,
x"000000E8" AFTER 11040 ns,
x"00000000" AFTER 11060 ns,
x"000000E4" AFTER 11080 ns,
x"00000000" AFTER 11100 ns,
x"000000E0" AFTER 11120 ns,
x"00000000" AFTER 11140 ns,
x"000000DC" AFTER 11160 ns,
x"00000000" AFTER 11180 ns,
x"000000D8" AFTER 11200 ns,
x"00000000" AFTER 11220 ns,
x"000000D4" AFTER 11240 ns,
x"00000000" AFTER 11260 ns,
x"000000D0" AFTER 11280 ns,
x"00000000" AFTER 11300 ns,
x"000000CC" AFTER 11320 ns,
x"00000000" AFTER 11340 ns,
x"000000C8" AFTER 11360 ns,
x"00000000" AFTER 11380 ns,
x"000000C4" AFTER 11400 ns,
x"00000000" AFTER 11420 ns,
x"000000C0" AFTER 11440 ns,
x"00000000" AFTER 11460 ns,
x"000000BC" AFTER 11480 ns,
x"00000000" AFTER 11500 ns,
x"000000B8" AFTER 11520 ns,
x"00000000" AFTER 11540 ns,
x"000000B4" AFTER 11560 ns,
x"00000000" AFTER 11580 ns,
x"000000B0" AFTER 11600 ns,
x"00000000" AFTER 11620 ns,
x"000000AC" AFTER 11640 ns,
x"00000000" AFTER 11660 ns,
x"000000A8" AFTER 11680 ns,
x"00000000" AFTER 11700 ns,
x"000000A4" AFTER 11720 ns,
x"00000000" AFTER 11740 ns,
x"000000A0" AFTER 11760 ns,
x"00000000" AFTER 11780 ns,
x"0000009C" AFTER 11800 ns,
x"00000000" AFTER 11820 ns,
x"00000098" AFTER 11840 ns,
x"00000000" AFTER 11860 ns,
x"00000094" AFTER 11880 ns,
x"00000000" AFTER 11900 ns,
x"00000090" AFTER 11920 ns,
x"00000000" AFTER 11940 ns,
x"0000008C" AFTER 11960 ns,
x"00000000" AFTER 11980 ns,
x"00000088" AFTER 12000 ns,
x"00000000" AFTER 12020 ns,
x"00000084" AFTER 12040 ns,
x"00000000" AFTER 12060 ns,
x"00000080" AFTER 12080 ns,
x"00000000" AFTER 12100 ns,
x"0000007C" AFTER 12120 ns,
x"00000000" AFTER 12140 ns,
x"00000078" AFTER 12160 ns,
x"00000000" AFTER 12180 ns,
x"00000074" AFTER 12200 ns,
x"00000000" AFTER 12220 ns,
x"00000070" AFTER 12240 ns,
x"00000000" AFTER 12260 ns,
x"0000006C" AFTER 12280 ns,
x"00000000" AFTER 12300 ns,
x"00000068" AFTER 12320 ns,
x"00000000" AFTER 12340 ns,
x"00000064" AFTER 12360 ns,
x"00000000" AFTER 12380 ns,
x"00000060" AFTER 12400 ns,
x"00000000" AFTER 12420 ns,
x"0000005C" AFTER 12440 ns,
x"00000000" AFTER 12460 ns,
x"00000058" AFTER 12480 ns,
x"00000000" AFTER 12500 ns,
x"00000054" AFTER 12520 ns,
x"00000000" AFTER 12540 ns,
x"00000050" AFTER 12560 ns,
x"00000000" AFTER 12580 ns,
x"0000004C" AFTER 12600 ns,
x"00000000" AFTER 12620 ns,
x"00000048" AFTER 12640 ns,
x"00000000" AFTER 12660 ns,
x"00000044" AFTER 12680 ns,
x"00000000" AFTER 12700 ns,
x"00000040" AFTER 12720 ns,
x"00000000" AFTER 12740 ns,
x"0000003C" AFTER 12760 ns,
x"00000000" AFTER 12780 ns,
x"00000038" AFTER 12800 ns,
x"00000000" AFTER 12820 ns,
x"00000034" AFTER 12840 ns,
x"00000000" AFTER 12860 ns,
x"00000030" AFTER 12880 ns,
x"00000000" AFTER 12900 ns,
x"0000002C" AFTER 12920 ns,
x"00000000" AFTER 12940 ns,
x"00000028" AFTER 12960 ns,
x"00000000" AFTER 12980 ns,
x"00000024" AFTER 13000 ns,
x"00000000" AFTER 13020 ns,
x"00000020" AFTER 13040 ns,
x"00000000" AFTER 13060 ns,
x"0000001C" AFTER 13080 ns,
x"00000000" AFTER 13100 ns,
x"00000018" AFTER 13120 ns,
x"00000000" AFTER 13140 ns,
x"00000014" AFTER 13160 ns,
x"00000000" AFTER 13180 ns,
x"00000010" AFTER 13200 ns,
x"00000000" AFTER 13220 ns,
x"0000000C" AFTER 13240 ns,
x"00000000" AFTER 13260 ns,
x"00000008" AFTER 13280 ns,
x"00000000" AFTER 13300 ns,
x"00000004" AFTER 13320 ns,
x"00000000" AFTER 13340 ns,
x"EE6B27FC" AFTER 13360 ns,
x"00000000" AFTER 13380 ns,
x"EE6B27F8" AFTER 13400 ns,
x"00000000" AFTER 13420 ns,
x"EE6B27F4" AFTER 13440 ns,
x"00000000" AFTER 13460 ns,
x"EE6B27F0" AFTER 13480 ns,
x"00000000" AFTER 13500 ns,
x"EE6B27EC" AFTER 13520 ns,
x"00000000" AFTER 13540 ns,
x"EE6B27E8" AFTER 13560 ns,
x"00000000" AFTER 13580 ns,
x"EE6B27E4" AFTER 13600 ns,
x"00000000" AFTER 13620 ns,
x"EE6B27E0" AFTER 13640 ns,
x"00000000" AFTER 13660 ns,
x"EE6B27DC" AFTER 13680 ns,
x"00000000" AFTER 13700 ns,
x"EE6B27D8" AFTER 13720 ns,
x"00000000" AFTER 13740 ns,
x"EE6B27D4" AFTER 13760 ns,
x"00000000" AFTER 13780 ns,
x"EE6B27D0" AFTER 13800 ns,
x"00000000" AFTER 13820 ns,
x"EE6B27CC" AFTER 13840 ns,
x"00000000" AFTER 13860 ns,
x"EE6B27C8" AFTER 13880 ns,
x"00000000" AFTER 13900 ns,
x"EE6B27C4" AFTER 13920 ns,
x"00000000" AFTER 13940 ns,
x"EE6B27C0" AFTER 13960 ns,
x"00000000" AFTER 13980 ns,
x"EE6B27BC" AFTER 14000 ns,
x"00000000" AFTER 14020 ns,
x"EE6B27B8" AFTER 14040 ns,
x"00000000" AFTER 14060 ns,
x"EE6B27B4" AFTER 14080 ns,
x"00000000" AFTER 14100 ns,
x"EE6B27B0" AFTER 14120 ns,
x"00000000" AFTER 14140 ns,
x"EE6B27AC" AFTER 14160 ns,
x"00000000" AFTER 14180 ns,
x"EE6B27A8" AFTER 14200 ns,
x"00000000" AFTER 14220 ns,
x"EE6B27A4" AFTER 14240 ns,
x"00000000" AFTER 14260 ns,
x"EE6B27A0" AFTER 14280 ns,
x"00000000" AFTER 14300 ns,
x"EE6B279C" AFTER 14320 ns,
x"00000000" AFTER 14340 ns,
x"EE6B2798" AFTER 14360 ns,
x"00000000" AFTER 14380 ns,
x"EE6B2794" AFTER 14400 ns,
x"00000000" AFTER 14420 ns,
x"EE6B2790" AFTER 14440 ns,
x"00000000" AFTER 14460 ns,
x"EE6B278C" AFTER 14480 ns,
x"00000000" AFTER 14500 ns,
x"EE6B2788" AFTER 14520 ns,
x"00000000" AFTER 14540 ns,
x"EE6B2784" AFTER 14560 ns,
x"00000000" AFTER 14580 ns,
x"EE6B2780" AFTER 14600 ns,
x"00000000" AFTER 14620 ns,
x"EE6B277C" AFTER 14640 ns,
x"00000000" AFTER 14660 ns,
x"EE6B2778" AFTER 14680 ns,
x"00000000" AFTER 14700 ns,
x"EE6B2774" AFTER 14720 ns,
x"00000000" AFTER 14740 ns,
x"EE6B2770" AFTER 14760 ns,
x"00000000" AFTER 14780 ns,
x"EE6B276C" AFTER 14800 ns,
x"00000000" AFTER 14820 ns,
x"EE6B2768" AFTER 14840 ns,
x"00000000" AFTER 14860 ns,
x"EE6B2764" AFTER 14880 ns,
x"00000000" AFTER 14900 ns,
x"EE6B2760" AFTER 14920 ns,
x"00000000" AFTER 14940 ns,
x"EE6B275C" AFTER 14960 ns,
x"00000000" AFTER 14980 ns,
x"EE6B2758" AFTER 15000 ns,
x"00000000" AFTER 15020 ns,
x"EE6B2754" AFTER 15040 ns,
x"00000000" AFTER 15060 ns,
x"EE6B2750" AFTER 15080 ns,
x"00000000" AFTER 15100 ns,
x"EE6B274C" AFTER 15120 ns,
x"00000000" AFTER 15140 ns,
x"EE6B2748" AFTER 15160 ns,
x"00000000" AFTER 15180 ns,
x"EE6B2744" AFTER 15200 ns,
x"00000000" AFTER 15220 ns,
x"EE6B2740" AFTER 15240 ns,
x"00000000" AFTER 15260 ns,
x"EE6B273C" AFTER 15280 ns,
x"00000000" AFTER 15300 ns,
x"EE6B2738" AFTER 15320 ns,
x"00000000" AFTER 15340 ns,
x"EE6B2734" AFTER 15360 ns,
x"00000000" AFTER 15380 ns,
x"EE6B2730" AFTER 15400 ns,
x"00000000" AFTER 15420 ns,
x"EE6B272C" AFTER 15440 ns,
x"00000000" AFTER 15460 ns,
x"EE6B2728" AFTER 15480 ns,
x"00000000" AFTER 15500 ns,
x"EE6B2724" AFTER 15520 ns,
x"00000000" AFTER 15540 ns,
x"EE6B2720" AFTER 15560 ns,
x"00000000" AFTER 15580 ns,
x"EE6B271C" AFTER 15600 ns,
x"00000000" AFTER 15620 ns,
x"EE6B2718" AFTER 15640 ns,
x"00000000" AFTER 15660 ns,
x"EE6B2714" AFTER 15680 ns,
x"00000000" AFTER 15700 ns,
x"EE6B2710" AFTER 15720 ns,
x"00000000" AFTER 15740 ns,
x"EE6B270C" AFTER 15760 ns,
x"00000000" AFTER 15780 ns,
x"EE6B2708" AFTER 15800 ns,
x"00000000" AFTER 15820 ns,
x"EE6B2704" AFTER 15840 ns,
x"00000000" AFTER 15860 ns,
x"EE6B2700" AFTER 15880 ns,
x"00000000" AFTER 15900 ns,
x"EE6B26FC" AFTER 15920 ns,
x"00000000" AFTER 15940 ns,
x"EE6B26F8" AFTER 15960 ns,
x"00000000" AFTER 15980 ns,
x"EE6B26F4" AFTER 16000 ns,
x"00000000" AFTER 16020 ns,
x"EE6B26F0" AFTER 16040 ns,
x"00000000" AFTER 16060 ns,
x"EE6B26EC" AFTER 16080 ns,
x"00000000" AFTER 16100 ns,
x"EE6B26E8" AFTER 16120 ns,
x"00000000" AFTER 16140 ns,
x"EE6B26E4" AFTER 16160 ns,
x"00000000" AFTER 16180 ns,
x"EE6B26E0" AFTER 16200 ns,
x"00000000" AFTER 16220 ns,
x"EE6B26DC" AFTER 16240 ns,
x"00000000" AFTER 16260 ns,
x"EE6B26D8" AFTER 16280 ns,
x"00000000" AFTER 16300 ns,
x"EE6B26D4" AFTER 16320 ns,
x"00000000" AFTER 16340 ns,
x"EE6B26D0" AFTER 16360 ns,
x"00000000" AFTER 16380 ns,
x"EE6B26CC" AFTER 16400 ns,
x"00000000" AFTER 16420 ns,
x"EE6B26C8" AFTER 16440 ns,
x"00000000" AFTER 16460 ns,
x"EE6B26C4" AFTER 16480 ns,
x"00000000" AFTER 16500 ns,
x"EE6B26C0" AFTER 16520 ns,
x"00000000" AFTER 16540 ns,
x"EE6B26BC" AFTER 16560 ns,
x"00000000" AFTER 16580 ns,
x"EE6B26B8" AFTER 16600 ns,
x"00000000" AFTER 16620 ns,
x"EE6B26B4" AFTER 16640 ns,
x"00000000" AFTER 16660 ns,
x"EE6B26B0" AFTER 16680 ns,
x"00000000" AFTER 16700 ns,
x"EE6B26AC" AFTER 16720 ns,
x"00000000" AFTER 16740 ns,
x"EE6B26A8" AFTER 16760 ns,
x"00000000" AFTER 16780 ns,
x"EE6B26A4" AFTER 16800 ns,
x"00000000" AFTER 16820 ns,
x"EE6B26A0" AFTER 16840 ns,
x"00000000" AFTER 16860 ns,
x"EE6B269C" AFTER 16880 ns,
x"00000000" AFTER 16900 ns,
x"EE6B2698" AFTER 16920 ns,
x"00000000" AFTER 16940 ns,
x"EE6B2694" AFTER 16960 ns,
x"00000000" AFTER 16980 ns,
x"EE6B2690" AFTER 17000 ns,
x"00000000" AFTER 17020 ns,
x"EE6B268C" AFTER 17040 ns,
x"00000000" AFTER 17060 ns,
x"EE6B2688" AFTER 17080 ns,
x"00000000" AFTER 17100 ns,
x"EE6B2684" AFTER 17120 ns,
x"00000000" AFTER 17140 ns,
x"EE6B2680" AFTER 17160 ns,
x"00000000" AFTER 17180 ns,
x"EE6B267C" AFTER 17200 ns,
x"00000000" AFTER 17220 ns,
x"EE6B2678" AFTER 17240 ns,
x"00000000" AFTER 17260 ns,
x"EE6B2674" AFTER 17280 ns,
x"00000000" AFTER 17300 ns,
x"EE6B2670" AFTER 17320 ns,
x"00000000" AFTER 17340 ns,
x"EE6B266C" AFTER 17360 ns,
x"00000000" AFTER 17380 ns,
x"EE6B2668" AFTER 17400 ns,
x"00000000" AFTER 17420 ns,
x"EE6B2664" AFTER 17440 ns,
x"00000000" AFTER 17460 ns,
x"EE6B2660" AFTER 17480 ns,
x"00000000" AFTER 17500 ns,
x"EE6B265C" AFTER 17520 ns,
x"00000000" AFTER 17540 ns,
x"EE6B2658" AFTER 17560 ns,
x"00000000" AFTER 17580 ns,
x"EE6B2654" AFTER 17600 ns,
x"00000000" AFTER 17620 ns,
x"EE6B2650" AFTER 17640 ns,
x"00000000" AFTER 17660 ns,
x"EE6B264C" AFTER 17680 ns,
x"00000000" AFTER 17700 ns,
x"EE6B2648" AFTER 17720 ns,
x"00000000" AFTER 17740 ns,
x"EE6B2644" AFTER 17760 ns,
x"00000000" AFTER 17780 ns,
x"EE6B2640" AFTER 17800 ns,
x"00000000" AFTER 17820 ns,
x"EE6B263C" AFTER 17840 ns,
x"00000000" AFTER 17860 ns,
x"EE6B2638" AFTER 17880 ns,
x"00000000" AFTER 17900 ns,
x"EE6B2634" AFTER 17920 ns,
x"00000000" AFTER 17940 ns,
x"EE6B2630" AFTER 17960 ns,
x"00000000" AFTER 17980 ns,
x"EE6B262C" AFTER 18000 ns,
x"00000000" AFTER 18020 ns,
x"EE6B2628" AFTER 18040 ns,
x"00000000" AFTER 18060 ns,
x"EE6B2624" AFTER 18080 ns,
x"00000000" AFTER 18100 ns,
x"EE6B2620" AFTER 18120 ns,
x"00000000" AFTER 18140 ns,
x"EE6B261C" AFTER 18160 ns,
x"00000000" AFTER 18180 ns,
x"EE6B2618" AFTER 18200 ns,
x"00000000" AFTER 18220 ns,
x"EE6B2614" AFTER 18240 ns,
x"00000000" AFTER 18260 ns,
x"EE6B2610" AFTER 18280 ns,
x"00000000" AFTER 18300 ns,
x"EE6B260C" AFTER 18320 ns,
x"00000000" AFTER 18340 ns,
x"EE6B2608" AFTER 18360 ns,
x"00000000" AFTER 18380 ns,
x"EE6B2604" AFTER 18400 ns,
x"00000000" AFTER 18420 ns,
x"EE6B2600" AFTER 18440 ns,
x"00000000" AFTER 18460 ns,
x"EE6B25FC" AFTER 18480 ns,
x"00000000" AFTER 18500 ns,
x"EE6B25F8" AFTER 18520 ns,
x"00000000" AFTER 18540 ns,
x"EE6B25F4" AFTER 18560 ns,
x"00000000" AFTER 18580 ns,
x"EE6B25F0" AFTER 18600 ns,
x"00000000" AFTER 18620 ns,
x"EE6B25EC" AFTER 18640 ns,
x"00000000" AFTER 18660 ns,
x"EE6B25E8" AFTER 18680 ns,
x"00000000" AFTER 18700 ns,
x"EE6B25E4" AFTER 18720 ns,
x"00000000" AFTER 18740 ns,
x"EE6B25E0" AFTER 18760 ns,
x"00000000" AFTER 18780 ns,
x"EE6B25DC" AFTER 18800 ns,
x"00000000" AFTER 18820 ns,
x"EE6B25D8" AFTER 18840 ns,
x"00000000" AFTER 18860 ns,
x"EE6B25D4" AFTER 18880 ns,
x"00000000" AFTER 18900 ns,
x"EE6B25D0" AFTER 18920 ns,
x"00000000" AFTER 18940 ns,
x"EE6B25CC" AFTER 18960 ns,
x"00000000" AFTER 18980 ns,
x"EE6B25C8" AFTER 19000 ns,
x"00000000" AFTER 19020 ns,
x"EE6B25C4" AFTER 19040 ns,
x"00000000" AFTER 19060 ns,
x"EE6B25C0" AFTER 19080 ns,
x"00000000" AFTER 19100 ns,
x"EE6B25BC" AFTER 19120 ns,
x"00000000" AFTER 19140 ns,
x"EE6B25B8" AFTER 19160 ns,
x"00000000" AFTER 19180 ns,
x"EE6B25B4" AFTER 19200 ns,
x"00000000" AFTER 19220 ns,
x"EE6B25B0" AFTER 19240 ns,
x"00000000" AFTER 19260 ns,
x"EE6B25AC" AFTER 19280 ns,
x"00000000" AFTER 19300 ns,
x"EE6B25A8" AFTER 19320 ns,
x"00000000" AFTER 19340 ns,
x"EE6B25A4" AFTER 19360 ns,
x"00000000" AFTER 19380 ns,
x"EE6B25A0" AFTER 19400 ns,
x"00000000" AFTER 19420 ns,
x"EE6B259C" AFTER 19440 ns,
x"00000000" AFTER 19460 ns,
x"EE6B2598" AFTER 19480 ns,
x"00000000" AFTER 19500 ns,
x"EE6B2594" AFTER 19520 ns,
x"00000000" AFTER 19540 ns,
x"EE6B2590" AFTER 19560 ns,
x"00000000" AFTER 19580 ns,
x"EE6B258C" AFTER 19600 ns,
x"00000000" AFTER 19620 ns,
x"EE6B2588" AFTER 19640 ns,
x"00000000" AFTER 19660 ns,
x"EE6B2584" AFTER 19680 ns,
x"00000000" AFTER 19700 ns,
x"EE6B2580" AFTER 19720 ns,
x"00000000" AFTER 19740 ns,
x"EE6B257C" AFTER 19760 ns,
x"00000000" AFTER 19780 ns,
x"EE6B2578" AFTER 19800 ns,
x"00000000" AFTER 19820 ns,
x"EE6B2574" AFTER 19840 ns,
x"00000000" AFTER 19860 ns,
x"EE6B2570" AFTER 19880 ns,
x"00000000" AFTER 19900 ns,
x"EE6B256C" AFTER 19920 ns,
x"00000000" AFTER 19940 ns,
x"EE6B2570" AFTER 19960 ns,
x"00000000" AFTER 19980 ns,
x"EE6B2574" AFTER 20000 ns,
x"00000000" AFTER 20020 ns,
x"EE6B2578" AFTER 20040 ns,
x"00000000" AFTER 20060 ns,
x"EE6B257C" AFTER 20080 ns,
x"00000000" AFTER 20100 ns,
x"EE6B2580" AFTER 20120 ns,
x"00000000" AFTER 20140 ns,
x"EE6B2584" AFTER 20160 ns,
x"00000000" AFTER 20180 ns,
x"EE6B2588" AFTER 20200 ns,
x"00000000" AFTER 20220 ns,
x"EE6B258C" AFTER 20240 ns,
x"00000000" AFTER 20260 ns,
x"EE6B2590" AFTER 20280 ns,
x"00000000" AFTER 20300 ns,
x"EE6B2594" AFTER 20320 ns,
x"00000000" AFTER 20340 ns,
x"EE6B2598" AFTER 20360 ns,
x"00000000" AFTER 20380 ns,
x"EE6B259C" AFTER 20400 ns,
x"00000000" AFTER 20420 ns,
x"EE6B25A0" AFTER 20440 ns,
x"00000000" AFTER 20460 ns,
x"EE6B25A4" AFTER 20480 ns,
x"00000000" AFTER 20500 ns,
x"EE6B25A8" AFTER 20520 ns,
x"00000000" AFTER 20540 ns,
x"EE6B25AC" AFTER 20560 ns,
x"00000000" AFTER 20580 ns,
x"EE6B25B0" AFTER 20600 ns,
x"00000000" AFTER 20620 ns,
x"EE6B25B4" AFTER 20640 ns,
x"00000000" AFTER 20660 ns,
x"EE6B25B8" AFTER 20680 ns,
x"00000000" AFTER 20700 ns,
x"EE6B25BC" AFTER 20720 ns,
x"00000000" AFTER 20740 ns,
x"EE6B25C0" AFTER 20760 ns,
x"00000000" AFTER 20780 ns,
x"EE6B25C4" AFTER 20800 ns,
x"00000000" AFTER 20820 ns,
x"EE6B25C8" AFTER 20840 ns,
x"00000000" AFTER 20860 ns,
x"EE6B25CC" AFTER 20880 ns,
x"00000000" AFTER 20900 ns,
x"EE6B25D0" AFTER 20920 ns,
x"00000000" AFTER 20940 ns,
x"EE6B25D4" AFTER 20960 ns,
x"00000000" AFTER 20980 ns,
x"EE6B25D8" AFTER 21000 ns,
x"00000000" AFTER 21020 ns,
x"EE6B25DC" AFTER 21040 ns,
x"00000000" AFTER 21060 ns,
x"EE6B25E0" AFTER 21080 ns,
x"00000000" AFTER 21100 ns,
x"EE6B25E4" AFTER 21120 ns,
x"00000000" AFTER 21140 ns,
x"EE6B25E8" AFTER 21160 ns,
x"00000000" AFTER 21180 ns,
x"EE6B25EC" AFTER 21200 ns,
x"00000000" AFTER 21220 ns,
x"EE6B25F0" AFTER 21240 ns,
x"00000000" AFTER 21260 ns,
x"EE6B25F4" AFTER 21280 ns,
x"00000000" AFTER 21300 ns,
x"EE6B25F8" AFTER 21320 ns,
x"00000000" AFTER 21340 ns,
x"EE6B25FC" AFTER 21360 ns,
x"00000000" AFTER 21380 ns,
x"EE6B2600" AFTER 21400 ns,
x"00000000" AFTER 21420 ns,
x"EE6B2604" AFTER 21440 ns,
x"00000000" AFTER 21460 ns,
x"EE6B2608" AFTER 21480 ns,
x"00000000" AFTER 21500 ns,
x"EE6B260C" AFTER 21520 ns,
x"00000000" AFTER 21540 ns,
x"EE6B2610" AFTER 21560 ns,
x"00000000" AFTER 21580 ns,
x"EE6B2614" AFTER 21600 ns,
x"00000000" AFTER 21620 ns,
x"EE6B2618" AFTER 21640 ns,
x"00000000" AFTER 21660 ns,
x"EE6B261C" AFTER 21680 ns,
x"00000000" AFTER 21700 ns,
x"EE6B2620" AFTER 21720 ns,
x"00000000" AFTER 21740 ns,
x"EE6B2624" AFTER 21760 ns,
x"00000000" AFTER 21780 ns,
x"EE6B2628" AFTER 21800 ns,
x"00000000" AFTER 21820 ns,
x"EE6B262C" AFTER 21840 ns,
x"00000000" AFTER 21860 ns,
x"EE6B2630" AFTER 21880 ns,
x"00000000" AFTER 21900 ns,
x"EE6B2634" AFTER 21920 ns,
x"00000000" AFTER 21940 ns,
x"EE6B2638" AFTER 21960 ns,
x"00000000" AFTER 21980 ns,
x"EE6B263C" AFTER 22000 ns,
x"00000000" AFTER 22020 ns,
x"EE6B2640" AFTER 22040 ns,
x"00000000" AFTER 22060 ns,
x"EE6B2644" AFTER 22080 ns,
x"00000000" AFTER 22100 ns,
x"EE6B2648" AFTER 22120 ns,
x"00000000" AFTER 22140 ns,
x"EE6B264C" AFTER 22160 ns,
x"00000000" AFTER 22180 ns,
x"EE6B2650" AFTER 22200 ns,
x"00000000" AFTER 22220 ns,
x"EE6B2654" AFTER 22240 ns,
x"00000000" AFTER 22260 ns,
x"EE6B2658" AFTER 22280 ns,
x"00000000" AFTER 22300 ns,
x"EE6B265C" AFTER 22320 ns,
x"00000000" AFTER 22340 ns,
x"EE6B2660" AFTER 22360 ns,
x"00000000" AFTER 22380 ns,
x"EE6B2664" AFTER 22400 ns,
x"00000000" AFTER 22420 ns,
x"EE6B2668" AFTER 22440 ns,
x"00000000" AFTER 22460 ns,
x"EE6B266C" AFTER 22480 ns,
x"00000000" AFTER 22500 ns,
x"EE6B2670" AFTER 22520 ns,
x"00000000" AFTER 22540 ns,
x"EE6B2674" AFTER 22560 ns,
x"00000000" AFTER 22580 ns,
x"EE6B2678" AFTER 22600 ns,
x"00000000" AFTER 22620 ns,
x"EE6B267C" AFTER 22640 ns,
x"00000000" AFTER 22660 ns,
x"EE6B2680" AFTER 22680 ns,
x"00000000" AFTER 22700 ns,
x"EE6B2684" AFTER 22720 ns,
x"00000000" AFTER 22740 ns,
x"EE6B2688" AFTER 22760 ns,
x"00000000" AFTER 22780 ns,
x"EE6B268C" AFTER 22800 ns,
x"00000000" AFTER 22820 ns,
x"EE6B2690" AFTER 22840 ns,
x"00000000" AFTER 22860 ns,
x"EE6B2694" AFTER 22880 ns,
x"00000000" AFTER 22900 ns,
x"EE6B2698" AFTER 22920 ns,
x"00000000" AFTER 22940 ns,
x"EE6B269C" AFTER 22960 ns,
x"00000000" AFTER 22980 ns,
x"EE6B26A0" AFTER 23000 ns,
x"00000000" AFTER 23020 ns,
x"EE6B26A4" AFTER 23040 ns,
x"00000000" AFTER 23060 ns,
x"EE6B26A8" AFTER 23080 ns,
x"00000000" AFTER 23100 ns,
x"EE6B26AC" AFTER 23120 ns,
x"00000000" AFTER 23140 ns,
x"EE6B26B0" AFTER 23160 ns,
x"00000000" AFTER 23180 ns,
x"EE6B26B4" AFTER 23200 ns,
x"00000000" AFTER 23220 ns,
x"EE6B26B8" AFTER 23240 ns,
x"00000000" AFTER 23260 ns,
x"EE6B26BC" AFTER 23280 ns,
x"00000000" AFTER 23300 ns,
x"EE6B26C0" AFTER 23320 ns,
x"00000000" AFTER 23340 ns,
x"EE6B26C4" AFTER 23360 ns,
x"00000000" AFTER 23380 ns,
x"EE6B26C8" AFTER 23400 ns,
x"00000000" AFTER 23420 ns,
x"EE6B26CC" AFTER 23440 ns,
x"00000000" AFTER 23460 ns,
x"EE6B26D0" AFTER 23480 ns,
x"00000000" AFTER 23500 ns,
x"EE6B26D4" AFTER 23520 ns,
x"00000000" AFTER 23540 ns,
x"EE6B26D8" AFTER 23560 ns,
x"00000000" AFTER 23580 ns,
x"EE6B26DC" AFTER 23600 ns,
x"00000000" AFTER 23620 ns,
x"EE6B26E0" AFTER 23640 ns,
x"00000000" AFTER 23660 ns,
x"EE6B26E4" AFTER 23680 ns,
x"00000000" AFTER 23700 ns,
x"EE6B26E8" AFTER 23720 ns,
x"00000000" AFTER 23740 ns,
x"EE6B26EC" AFTER 23760 ns,
x"00000000" AFTER 23780 ns,
x"EE6B26F0" AFTER 23800 ns,
x"00000000" AFTER 23820 ns,
x"EE6B26F4" AFTER 23840 ns,
x"00000000" AFTER 23860 ns,
x"EE6B26F8" AFTER 23880 ns,
x"00000000" AFTER 23900 ns,
x"EE6B26FC" AFTER 23920 ns,
x"00000000" AFTER 23940 ns,
x"EE6B2700" AFTER 23960 ns,
x"00000000" AFTER 23980 ns,
x"EE6B2704" AFTER 24000 ns,
x"00000000" AFTER 24020 ns,
x"EE6B2708" AFTER 24040 ns,
x"00000000" AFTER 24060 ns,
x"EE6B270C" AFTER 24080 ns,
x"00000000" AFTER 24100 ns,
x"EE6B2710" AFTER 24120 ns,
x"00000000" AFTER 24140 ns,
x"EE6B2714" AFTER 24160 ns,
x"00000000" AFTER 24180 ns,
x"EE6B2718" AFTER 24200 ns,
x"00000000" AFTER 24220 ns,
x"EE6B271C" AFTER 24240 ns,
x"00000000" AFTER 24260 ns,
x"EE6B2720" AFTER 24280 ns,
x"00000000" AFTER 24300 ns,
x"EE6B2724" AFTER 24320 ns,
x"00000000" AFTER 24340 ns,
x"EE6B2728" AFTER 24360 ns,
x"00000000" AFTER 24380 ns,
x"EE6B272C" AFTER 24400 ns,
x"00000000" AFTER 24420 ns,
x"EE6B2730" AFTER 24440 ns,
x"00000000" AFTER 24460 ns,
x"EE6B2734" AFTER 24480 ns,
x"00000000" AFTER 24500 ns,
x"EE6B2738" AFTER 24520 ns,
x"00000000" AFTER 24540 ns,
x"EE6B273C" AFTER 24560 ns,
x"00000000" AFTER 24580 ns,
x"EE6B2740" AFTER 24600 ns,
x"00000000" AFTER 24620 ns,
x"EE6B2744" AFTER 24640 ns,
x"00000000" AFTER 24660 ns,
x"EE6B2748" AFTER 24680 ns,
x"00000000" AFTER 24700 ns,
x"EE6B274C" AFTER 24720 ns,
x"00000000" AFTER 24740 ns,
x"EE6B2750" AFTER 24760 ns,
x"00000000" AFTER 24780 ns,
x"EE6B2754" AFTER 24800 ns,
x"00000000" AFTER 24820 ns,
x"EE6B2758" AFTER 24840 ns,
x"00000000" AFTER 24860 ns,
x"EE6B275C" AFTER 24880 ns,
x"00000000" AFTER 24900 ns,
x"EE6B2760" AFTER 24920 ns,
x"00000000" AFTER 24940 ns,
x"EE6B2764" AFTER 24960 ns,
x"00000000" AFTER 24980 ns,
x"EE6B2768" AFTER 25000 ns,
x"00000000" AFTER 25020 ns,
x"EE6B276C" AFTER 25040 ns,
x"00000000" AFTER 25060 ns,
x"EE6B2770" AFTER 25080 ns,
x"00000000" AFTER 25100 ns,
x"EE6B2774" AFTER 25120 ns,
x"00000000" AFTER 25140 ns,
x"EE6B2778" AFTER 25160 ns,
x"00000000" AFTER 25180 ns,
x"EE6B277C" AFTER 25200 ns,
x"00000000" AFTER 25220 ns,
x"EE6B2780" AFTER 25240 ns,
x"00000000" AFTER 25260 ns,
x"EE6B2784" AFTER 25280 ns,
x"00000000" AFTER 25300 ns,
x"EE6B2788" AFTER 25320 ns,
x"00000000" AFTER 25340 ns,
x"EE6B278C" AFTER 25360 ns,
x"00000000" AFTER 25380 ns,
x"EE6B2790" AFTER 25400 ns,
x"00000000" AFTER 25420 ns,
x"EE6B2794" AFTER 25440 ns,
x"00000000" AFTER 25460 ns,
x"EE6B2798" AFTER 25480 ns,
x"00000000" AFTER 25500 ns,
x"EE6B279C" AFTER 25520 ns,
x"00000000" AFTER 25540 ns,
x"EE6B27A0" AFTER 25560 ns,
x"00000000" AFTER 25580 ns,
x"EE6B27A4" AFTER 25600 ns,
x"00000000" AFTER 25620 ns,
x"EE6B27A8" AFTER 25640 ns,
x"00000000" AFTER 25660 ns,
x"EE6B27AC" AFTER 25680 ns,
x"00000000" AFTER 25700 ns,
x"EE6B27B0" AFTER 25720 ns,
x"00000000" AFTER 25740 ns,
x"EE6B27B4" AFTER 25760 ns,
x"00000000" AFTER 25780 ns,
x"EE6B27B8" AFTER 25800 ns,
x"00000000" AFTER 25820 ns,
x"EE6B27BC" AFTER 25840 ns,
x"00000000" AFTER 25860 ns,
x"EE6B27C0" AFTER 25880 ns,
x"00000000" AFTER 25900 ns,
x"EE6B27C4" AFTER 25920 ns,
x"00000000" AFTER 25940 ns,
x"EE6B27C8" AFTER 25960 ns,
x"00000000" AFTER 25980 ns,
x"EE6B27CC" AFTER 26000 ns,
x"00000000" AFTER 26020 ns,
x"EE6B27D0" AFTER 26040 ns,
x"00000000" AFTER 26060 ns,
x"EE6B27D4" AFTER 26080 ns,
x"00000000" AFTER 26100 ns,
x"EE6B27D8" AFTER 26120 ns,
x"00000000" AFTER 26140 ns,
x"EE6B27DC" AFTER 26160 ns,
x"00000000" AFTER 26180 ns,
x"EE6B27E0" AFTER 26200 ns,
x"00000000" AFTER 26220 ns,
x"EE6B27E4" AFTER 26240 ns,
x"00000000" AFTER 26260 ns,
x"EE6B27E8" AFTER 26280 ns,
x"00000000" AFTER 26300 ns,
x"EE6B27EC" AFTER 26320 ns,
x"00000000" AFTER 26340 ns,
x"EE6B27F0" AFTER 26360 ns,
x"00000000" AFTER 26380 ns,
x"EE6B27F4" AFTER 26400 ns,
x"00000000" AFTER 26420 ns,
x"EE6B27F8" AFTER 26440 ns,
x"00000000" AFTER 26460 ns,
x"EE6B27FC" AFTER 26480 ns,
x"00000000" AFTER 26500 ns,
x"EE6B2800" AFTER 26520 ns,
x"00000000" AFTER 26540 ns,
x"EE6B2804" AFTER 26560 ns,
x"00000000" AFTER 26580 ns,
x"EE6B2808" AFTER 26600 ns,
x"00000000" AFTER 26620 ns,
x"EE6B280C" AFTER 26640 ns,
x"00000000" AFTER 26660 ns,
x"EE6B2810" AFTER 26680 ns,
x"00000000" AFTER 26700 ns,
x"EE6B2814" AFTER 26720 ns,
x"00000000" AFTER 26740 ns,
x"EE6B2818" AFTER 26760 ns,
x"00000000" AFTER 26780 ns,
x"EE6B281C" AFTER 26800 ns,
x"00000000" AFTER 26820 ns,
x"EE6B2820" AFTER 26840 ns,
x"00000000" AFTER 26860 ns,
x"EE6B2824" AFTER 26880 ns,
x"00000000" AFTER 26900 ns,
x"EE6B2828" AFTER 26920 ns,
x"00000000" AFTER 26940 ns,
x"EE6B282C" AFTER 26960 ns,
x"00000000" AFTER 26980 ns,
x"EE6B2830" AFTER 27000 ns,
x"00000000" AFTER 27020 ns,
x"EE6B2834" AFTER 27040 ns,
x"00000000" AFTER 27060 ns,
x"EE6B2838" AFTER 27080 ns,
x"00000000" AFTER 27100 ns,
x"EE6B283C" AFTER 27120 ns,
x"00000000" AFTER 27140 ns,
x"EE6B2840" AFTER 27160 ns,
x"00000000" AFTER 27180 ns,
x"EE6B2844" AFTER 27200 ns,
x"00000000" AFTER 27220 ns,
x"EE6B2848" AFTER 27240 ns,
x"00000000" AFTER 27260 ns,
x"EE6B284C" AFTER 27280 ns,
x"00000000" AFTER 27300 ns,
x"EE6B2850" AFTER 27320 ns,
x"00000000" AFTER 27340 ns,
x"EE6B2854" AFTER 27360 ns,
x"00000000" AFTER 27380 ns,
x"EE6B2858" AFTER 27400 ns,
x"00000000" AFTER 27420 ns,
x"EE6B285C" AFTER 27440 ns,
x"00000000" AFTER 27460 ns,
x"EE6B2860" AFTER 27480 ns,
x"00000000" AFTER 27500 ns,
x"EE6B2864" AFTER 27520 ns,
x"00000000" AFTER 27540 ns,
x"EE6B2868" AFTER 27560 ns,
x"00000000" AFTER 27580 ns,
x"EE6B286C" AFTER 27600 ns,
x"00000000" AFTER 27620 ns,
x"EE6B2870" AFTER 27640 ns,
x"00000000" AFTER 27660 ns,
x"EE6B2874" AFTER 27680 ns,
x"00000000" AFTER 27700 ns,
x"EE6B2878" AFTER 27720 ns,
x"00000000" AFTER 27740 ns,
x"EE6B287C" AFTER 27760 ns,
x"00000000" AFTER 27780 ns,
x"EE6B2880" AFTER 27800 ns,
x"00000000" AFTER 27820 ns,
x"EE6B2884" AFTER 27840 ns,
x"00000000" AFTER 27860 ns,
x"EE6B2888" AFTER 27880 ns,
x"00000000" AFTER 27900 ns,
x"EE6B288C" AFTER 27920 ns,
x"00000000" AFTER 27940 ns,
x"EE6B2890" AFTER 27960 ns,
x"00000000" AFTER 27980 ns,
x"EE6B2894" AFTER 28000 ns,
x"00000000" AFTER 28020 ns,
x"EE6B2898" AFTER 28040 ns,
x"00000000" AFTER 28060 ns,
x"EE6B289C" AFTER 28080 ns,
x"00000000" AFTER 28100 ns,
x"EE6B28A0" AFTER 28120 ns,
x"00000000" AFTER 28140 ns,
x"EE6B28A4" AFTER 28160 ns,
x"00000000" AFTER 28180 ns,
x"EE6B28A8" AFTER 28200 ns,
x"00000000" AFTER 28220 ns,
x"EE6B28AC" AFTER 28240 ns,
x"00000000" AFTER 28260 ns,
x"EE6B28B0" AFTER 28280 ns,
x"00000000" AFTER 28300 ns,
x"EE6B28B4" AFTER 28320 ns,
x"00000000" AFTER 28340 ns,
x"EE6B28B8" AFTER 28360 ns,
x"00000000" AFTER 28380 ns,
x"EE6B28BC" AFTER 28400 ns,
x"00000000" AFTER 28420 ns,
x"EE6B28C0" AFTER 28440 ns,
x"00000000" AFTER 28460 ns,
x"EE6B28C4" AFTER 28480 ns,
x"00000000" AFTER 28500 ns,
x"EE6B28C8" AFTER 28520 ns,
x"00000000" AFTER 28540 ns,
x"EE6B28CC" AFTER 28560 ns,
x"00000000" AFTER 28580 ns,
x"EE6B28D0" AFTER 28600 ns,
x"00000000" AFTER 28620 ns,
x"EE6B28D4" AFTER 28640 ns,
x"00000000" AFTER 28660 ns,
x"EE6B28D8" AFTER 28680 ns,
x"00000000" AFTER 28700 ns,
x"EE6B28DC" AFTER 28720 ns,
x"00000000" AFTER 28740 ns,
x"EE6B28E0" AFTER 28760 ns,
x"00000000" AFTER 28780 ns,
x"EE6B28E4" AFTER 28800 ns,
x"00000000" AFTER 28820 ns,
x"EE6B28E8" AFTER 28840 ns,
x"00000000" AFTER 28860 ns,
x"EE6B28EC" AFTER 28880 ns,
x"00000000" AFTER 28900 ns,
x"EE6B28F0" AFTER 28920 ns,
x"00000000" AFTER 28940 ns,
x"EE6B28F4" AFTER 28960 ns,
x"00000000" AFTER 28980 ns,
x"EE6B28F8" AFTER 29000 ns,
x"00000000" AFTER 29020 ns,
x"EE6B28FC" AFTER 29040 ns,
x"00000000" AFTER 29060 ns,
x"EE6B2900" AFTER 29080 ns,
x"00000000" AFTER 29100 ns,
x"EE6B2904" AFTER 29120 ns,
x"00000000" AFTER 29140 ns,
x"EE6B2908" AFTER 29160 ns,
x"00000000" AFTER 29180 ns,
x"EE6B290C" AFTER 29200 ns,
x"00000000" AFTER 29220 ns,
x"EE6B2910" AFTER 29240 ns,
x"00000000" AFTER 29260 ns,
x"EE6B2914" AFTER 29280 ns,
x"00000000" AFTER 29300 ns,
x"EE6B2918" AFTER 29320 ns,
x"00000000" AFTER 29340 ns,
x"EE6B291C" AFTER 29360 ns,
x"00000000" AFTER 29380 ns,
x"EE6B2920" AFTER 29400 ns,
x"00000000" AFTER 29420 ns,
x"EE6B2924" AFTER 29440 ns,
x"00000000" AFTER 29460 ns,
x"EE6B2928" AFTER 29480 ns,
x"00000000" AFTER 29500 ns,
x"EE6B292C" AFTER 29520 ns,
x"00000000" AFTER 29540 ns,
x"EE6B2930" AFTER 29560 ns,
x"00000000" AFTER 29580 ns,
x"EE6B2934" AFTER 29600 ns,
x"00000000" AFTER 29620 ns,
x"EE6B2938" AFTER 29640 ns,
x"00000000" AFTER 29660 ns,
x"EE6B293C" AFTER 29680 ns,
x"00000000" AFTER 29700 ns,
x"EE6B2940" AFTER 29720 ns,
x"00000000" AFTER 29740 ns,
x"EE6B2944" AFTER 29760 ns,
x"00000000" AFTER 29780 ns,
x"EE6B2948" AFTER 29800 ns,
x"00000000" AFTER 29820 ns,
x"EE6B294C" AFTER 29840 ns,
x"00000000" AFTER 29860 ns,
x"EE6B2950" AFTER 29880 ns,
x"00000000" AFTER 29900 ns,
x"EE6B2954" AFTER 29920 ns,
x"00000000" AFTER 29940 ns,
x"EE6B2958" AFTER 29960 ns,
x"00000000" AFTER 29980 ns,
x"EE6B295C" AFTER 30000 ns,
x"00000000" AFTER 30020 ns,
x"EE6B2960" AFTER 30040 ns,
x"00000000" AFTER 30060 ns,
x"EE6B2964" AFTER 30080 ns,
x"00000000" AFTER 30100 ns,
x"EE6B2968" AFTER 30120 ns,
x"00000000" AFTER 30140 ns,
x"EE6B296C" AFTER 30160 ns,
x"00000000" AFTER 30180 ns,
x"EE6B2970" AFTER 30200 ns,
x"00000000" AFTER 30220 ns,
x"EE6B2974" AFTER 30240 ns,
x"00000000" AFTER 30260 ns,
x"EE6B2978" AFTER 30280 ns,
x"00000000" AFTER 30300 ns,
x"EE6B297C" AFTER 30320 ns,
x"00000000" AFTER 30340 ns,
x"EE6B2980" AFTER 30360 ns,
x"00000000" AFTER 30380 ns,
x"EE6B2984" AFTER 30400 ns,
x"00000000" AFTER 30420 ns,
x"EE6B2988" AFTER 30440 ns,
x"00000000" AFTER 30460 ns,
x"EE6B298C" AFTER 30480 ns,
x"00000000" AFTER 30500 ns,
x"EE6B2990" AFTER 30520 ns,
x"00000000" AFTER 30540 ns,
x"EE6B2994" AFTER 30560 ns,
x"00000000" AFTER 30580 ns,
x"EE6B2998" AFTER 30600 ns,
x"00000000" AFTER 30620 ns,
x"EE6B299C" AFTER 30640 ns,
x"00000000" AFTER 30660 ns,
x"EE6B29A0" AFTER 30680 ns,
x"00000000" AFTER 30700 ns,
x"EE6B29A4" AFTER 30720 ns,
x"00000000" AFTER 30740 ns,
x"EE6B29A8" AFTER 30760 ns,
x"00000000" AFTER 30780 ns,
x"EE6B29AC" AFTER 30800 ns,
x"00000000" AFTER 30820 ns,
x"EE6B29B0" AFTER 30840 ns,
x"00000000" AFTER 30860 ns,
x"EE6B29B4" AFTER 30880 ns,
x"00000000" AFTER 30900 ns,
x"EE6B29B8" AFTER 30920 ns,
x"00000000" AFTER 30940 ns,
x"EE6B29BC" AFTER 30960 ns;

AluRegisters <= x"00000000" AFTER 00020 ns,
x"00000532" AFTER 00040 ns,
x"00000000" AFTER 00060 ns,
x"0000052E" AFTER 00080 ns,
x"00000000" AFTER 00100 ns,
x"0000052A" AFTER 00120 ns,
x"00000000" AFTER 00140 ns,
x"00000526" AFTER 00160 ns,
x"00000000" AFTER 00180 ns,
x"00000522" AFTER 00200 ns,
x"00000000" AFTER 00220 ns,
x"0000051E" AFTER 00240 ns,
x"00000000" AFTER 00260 ns,
x"0000051A" AFTER 00280 ns,
x"00000000" AFTER 00300 ns,
x"00000516" AFTER 00320 ns,
x"00000000" AFTER 00340 ns,
x"00000512" AFTER 00360 ns,
x"00000000" AFTER 00380 ns,
x"0000050E" AFTER 00400 ns,
x"00000000" AFTER 00420 ns,
x"0000050A" AFTER 00440 ns,
x"00000000" AFTER 00460 ns,
x"00000506" AFTER 00480 ns,
x"00000000" AFTER 00500 ns,
x"00000502" AFTER 00520 ns,
x"00000000" AFTER 00540 ns,
x"000004FE" AFTER 00560 ns,
x"00000000" AFTER 00580 ns,
x"000004FA" AFTER 00600 ns,
x"00000000" AFTER 00620 ns,
x"000004F6" AFTER 00640 ns,
x"00000000" AFTER 00660 ns,
x"000004F2" AFTER 00680 ns,
x"00000000" AFTER 00700 ns,
x"000004EE" AFTER 00720 ns,
x"00000000" AFTER 00740 ns,
x"000004EA" AFTER 00760 ns,
x"00000000" AFTER 00780 ns,
x"000004E6" AFTER 00800 ns,
x"00000000" AFTER 00820 ns,
x"000004E2" AFTER 00840 ns,
x"00000000" AFTER 00860 ns,
x"000004DE" AFTER 00880 ns,
x"00000000" AFTER 00900 ns,
x"000004DA" AFTER 00920 ns,
x"00000000" AFTER 00940 ns,
x"000004D6" AFTER 00960 ns,
x"00000000" AFTER 00980 ns,
x"000004D2" AFTER 01000 ns,
x"00000000" AFTER 01020 ns,
x"000004CE" AFTER 01040 ns,
x"00000000" AFTER 01060 ns,
x"000004CA" AFTER 01080 ns,
x"00000000" AFTER 01100 ns,
x"000004C6" AFTER 01120 ns,
x"00000000" AFTER 01140 ns,
x"000004C2" AFTER 01160 ns,
x"00000000" AFTER 01180 ns,
x"000004BE" AFTER 01200 ns,
x"00000000" AFTER 01220 ns,
x"000004BA" AFTER 01240 ns,
x"00000000" AFTER 01260 ns,
x"000004B6" AFTER 01280 ns,
x"00000000" AFTER 01300 ns,
x"000004B2" AFTER 01320 ns,
x"00000000" AFTER 01340 ns,
x"000004AE" AFTER 01360 ns,
x"00000000" AFTER 01380 ns,
x"000004AA" AFTER 01400 ns,
x"00000000" AFTER 01420 ns,
x"000004A6" AFTER 01440 ns,
x"00000000" AFTER 01460 ns,
x"000004A2" AFTER 01480 ns,
x"00000000" AFTER 01500 ns,
x"0000049E" AFTER 01520 ns,
x"00000000" AFTER 01540 ns,
x"0000049A" AFTER 01560 ns,
x"00000000" AFTER 01580 ns,
x"00000496" AFTER 01600 ns,
x"00000000" AFTER 01620 ns,
x"00000492" AFTER 01640 ns,
x"00000000" AFTER 01660 ns,
x"0000048E" AFTER 01680 ns,
x"00000000" AFTER 01700 ns,
x"0000048A" AFTER 01720 ns,
x"00000000" AFTER 01740 ns,
x"00000486" AFTER 01760 ns,
x"00000000" AFTER 01780 ns,
x"00000482" AFTER 01800 ns,
x"00000000" AFTER 01820 ns,
x"0000047E" AFTER 01840 ns,
x"00000000" AFTER 01860 ns,
x"0000047A" AFTER 01880 ns,
x"00000000" AFTER 01900 ns,
x"00000476" AFTER 01920 ns,
x"00000000" AFTER 01940 ns,
x"00000472" AFTER 01960 ns,
x"00000000" AFTER 01980 ns,
x"0000046E" AFTER 02000 ns,
x"00000000" AFTER 02020 ns,
x"0000046A" AFTER 02040 ns,
x"00000000" AFTER 02060 ns,
x"00000466" AFTER 02080 ns,
x"00000000" AFTER 02100 ns,
x"00000462" AFTER 02120 ns,
x"00000000" AFTER 02140 ns,
x"0000045E" AFTER 02160 ns,
x"00000000" AFTER 02180 ns,
x"0000045A" AFTER 02200 ns,
x"00000000" AFTER 02220 ns,
x"00000456" AFTER 02240 ns,
x"00000000" AFTER 02260 ns,
x"00000452" AFTER 02280 ns,
x"00000000" AFTER 02300 ns,
x"0000044E" AFTER 02320 ns,
x"00000000" AFTER 02340 ns,
x"0000044A" AFTER 02360 ns,
x"00000000" AFTER 02380 ns,
x"00000446" AFTER 02400 ns,
x"00000000" AFTER 02420 ns,
x"00000442" AFTER 02440 ns,
x"00000000" AFTER 02460 ns,
x"0000043E" AFTER 02480 ns,
x"00000000" AFTER 02500 ns,
x"0000043A" AFTER 02520 ns,
x"00000000" AFTER 02540 ns,
x"00000436" AFTER 02560 ns,
x"00000000" AFTER 02580 ns,
x"00000432" AFTER 02600 ns,
x"00000000" AFTER 02620 ns,
x"0000042E" AFTER 02640 ns,
x"00000000" AFTER 02660 ns,
x"0000042A" AFTER 02680 ns,
x"00000000" AFTER 02700 ns,
x"00000426" AFTER 02720 ns,
x"00000000" AFTER 02740 ns,
x"00000422" AFTER 02760 ns,
x"00000000" AFTER 02780 ns,
x"0000041E" AFTER 02800 ns,
x"00000000" AFTER 02820 ns,
x"0000041A" AFTER 02840 ns,
x"00000000" AFTER 02860 ns,
x"00000416" AFTER 02880 ns,
x"00000000" AFTER 02900 ns,
x"00000412" AFTER 02920 ns,
x"00000000" AFTER 02940 ns,
x"0000040E" AFTER 02960 ns,
x"00000000" AFTER 02980 ns,
x"0000040A" AFTER 03000 ns,
x"00000000" AFTER 03020 ns,
x"00000406" AFTER 03040 ns,
x"00000000" AFTER 03060 ns,
x"00000402" AFTER 03080 ns,
x"00000000" AFTER 03100 ns,
x"000003FE" AFTER 03120 ns,
x"00000000" AFTER 03140 ns,
x"000003FA" AFTER 03160 ns,
x"00000000" AFTER 03180 ns,
x"000003F6" AFTER 03200 ns,
x"00000000" AFTER 03220 ns,
x"000003F2" AFTER 03240 ns,
x"00000000" AFTER 03260 ns,
x"000003EE" AFTER 03280 ns,
x"00000000" AFTER 03300 ns,
x"000003EA" AFTER 03320 ns,
x"00000000" AFTER 03340 ns,
x"000003E6" AFTER 03360 ns,
x"00000000" AFTER 03380 ns,
x"000003E2" AFTER 03400 ns,
x"00000000" AFTER 03420 ns,
x"000003DE" AFTER 03440 ns,
x"00000000" AFTER 03460 ns,
x"000003DA" AFTER 03480 ns,
x"00000000" AFTER 03500 ns,
x"000003D6" AFTER 03520 ns,
x"00000000" AFTER 03540 ns,
x"000003D2" AFTER 03560 ns,
x"00000000" AFTER 03580 ns,
x"000003CE" AFTER 03600 ns,
x"00000000" AFTER 03620 ns,
x"000003CA" AFTER 03640 ns,
x"00000000" AFTER 03660 ns,
x"000003C6" AFTER 03680 ns,
x"00000000" AFTER 03700 ns,
x"000003C2" AFTER 03720 ns,
x"00000000" AFTER 03740 ns,
x"000003BE" AFTER 03760 ns,
x"00000000" AFTER 03780 ns,
x"000003BA" AFTER 03800 ns,
x"00000000" AFTER 03820 ns,
x"000003B6" AFTER 03840 ns,
x"00000000" AFTER 03860 ns,
x"000003B2" AFTER 03880 ns,
x"00000000" AFTER 03900 ns,
x"000003AE" AFTER 03920 ns,
x"00000000" AFTER 03940 ns,
x"000003AA" AFTER 03960 ns,
x"00000000" AFTER 03980 ns,
x"000003A6" AFTER 04000 ns,
x"00000000" AFTER 04020 ns,
x"000003A2" AFTER 04040 ns,
x"00000000" AFTER 04060 ns,
x"0000039E" AFTER 04080 ns,
x"00000000" AFTER 04100 ns,
x"0000039A" AFTER 04120 ns,
x"00000000" AFTER 04140 ns,
x"00000396" AFTER 04160 ns,
x"00000000" AFTER 04180 ns,
x"00000392" AFTER 04200 ns,
x"00000000" AFTER 04220 ns,
x"0000038E" AFTER 04240 ns,
x"00000000" AFTER 04260 ns,
x"0000038A" AFTER 04280 ns,
x"00000000" AFTER 04300 ns,
x"00000386" AFTER 04320 ns,
x"00000000" AFTER 04340 ns,
x"00000382" AFTER 04360 ns,
x"00000000" AFTER 04380 ns,
x"0000037E" AFTER 04400 ns,
x"00000000" AFTER 04420 ns,
x"0000037A" AFTER 04440 ns,
x"00000000" AFTER 04460 ns,
x"00000376" AFTER 04480 ns,
x"00000000" AFTER 04500 ns,
x"00000372" AFTER 04520 ns,
x"00000000" AFTER 04540 ns,
x"0000036E" AFTER 04560 ns,
x"00000000" AFTER 04580 ns,
x"0000036A" AFTER 04600 ns,
x"00000000" AFTER 04620 ns,
x"00000366" AFTER 04640 ns,
x"00000000" AFTER 04660 ns,
x"00000362" AFTER 04680 ns,
x"00000000" AFTER 04700 ns,
x"0000035E" AFTER 04720 ns,
x"00000000" AFTER 04740 ns,
x"0000035A" AFTER 04760 ns,
x"00000000" AFTER 04780 ns,
x"00000356" AFTER 04800 ns,
x"00000000" AFTER 04820 ns,
x"00000352" AFTER 04840 ns,
x"00000000" AFTER 04860 ns,
x"0000034E" AFTER 04880 ns,
x"00000000" AFTER 04900 ns,
x"0000034A" AFTER 04920 ns,
x"00000000" AFTER 04940 ns,
x"00000346" AFTER 04960 ns,
x"00000000" AFTER 04980 ns,
x"00000342" AFTER 05000 ns,
x"00000000" AFTER 05020 ns,
x"0000033E" AFTER 05040 ns,
x"00000000" AFTER 05060 ns,
x"0000033A" AFTER 05080 ns,
x"00000000" AFTER 05100 ns,
x"00000336" AFTER 05120 ns,
x"00000000" AFTER 05140 ns,
x"00000332" AFTER 05160 ns,
x"00000000" AFTER 05180 ns,
x"0000032E" AFTER 05200 ns,
x"00000000" AFTER 05220 ns,
x"0000032A" AFTER 05240 ns,
x"00000000" AFTER 05260 ns,
x"00000326" AFTER 05280 ns,
x"00000000" AFTER 05300 ns,
x"00000322" AFTER 05320 ns,
x"00000000" AFTER 05340 ns,
x"0000031E" AFTER 05360 ns,
x"00000000" AFTER 05380 ns,
x"0000031A" AFTER 05400 ns,
x"00000000" AFTER 05420 ns,
x"00000316" AFTER 05440 ns,
x"00000000" AFTER 05460 ns,
x"00000312" AFTER 05480 ns,
x"00000000" AFTER 05500 ns,
x"0000030E" AFTER 05520 ns,
x"00000000" AFTER 05540 ns,
x"0000030A" AFTER 05560 ns,
x"00000000" AFTER 05580 ns,
x"00000306" AFTER 05600 ns,
x"00000000" AFTER 05620 ns,
x"00000302" AFTER 05640 ns,
x"00000000" AFTER 05660 ns,
x"000002FE" AFTER 05680 ns,
x"00000000" AFTER 05700 ns,
x"000002FA" AFTER 05720 ns,
x"00000000" AFTER 05740 ns,
x"000002F6" AFTER 05760 ns,
x"00000000" AFTER 05780 ns,
x"000002F2" AFTER 05800 ns,
x"00000000" AFTER 05820 ns,
x"000002EE" AFTER 05840 ns,
x"00000000" AFTER 05860 ns,
x"000002EA" AFTER 05880 ns,
x"00000000" AFTER 05900 ns,
x"000002E6" AFTER 05920 ns,
x"00000000" AFTER 05940 ns,
x"000002E2" AFTER 05960 ns,
x"00000000" AFTER 05980 ns,
x"000002DE" AFTER 06000 ns,
x"00000000" AFTER 06020 ns,
x"000002DA" AFTER 06040 ns,
x"00000000" AFTER 06060 ns,
x"000002D6" AFTER 06080 ns,
x"00000000" AFTER 06100 ns,
x"000002D2" AFTER 06120 ns,
x"00000000" AFTER 06140 ns,
x"000002CE" AFTER 06160 ns,
x"00000000" AFTER 06180 ns,
x"000002CA" AFTER 06200 ns,
x"00000000" AFTER 06220 ns,
x"000002C6" AFTER 06240 ns,
x"00000000" AFTER 06260 ns,
x"000002C2" AFTER 06280 ns,
x"00000000" AFTER 06300 ns,
x"000002BE" AFTER 06320 ns,
x"00000000" AFTER 06340 ns,
x"000002BA" AFTER 06360 ns,
x"00000000" AFTER 06380 ns,
x"000002B6" AFTER 06400 ns,
x"00000000" AFTER 06420 ns,
x"000002B2" AFTER 06440 ns,
x"00000000" AFTER 06460 ns,
x"000002AE" AFTER 06480 ns,
x"00000000" AFTER 06500 ns,
x"000002AA" AFTER 06520 ns,
x"00000000" AFTER 06540 ns,
x"000002A6" AFTER 06560 ns,
x"00000000" AFTER 06580 ns,
x"000002A2" AFTER 06600 ns,
x"00000000" AFTER 06620 ns,
x"0000029E" AFTER 06640 ns,
x"00000000" AFTER 06660 ns,
x"0000029A" AFTER 06680 ns,
x"00000000" AFTER 06700 ns,
x"00000296" AFTER 06720 ns,
x"00000000" AFTER 06740 ns,
x"00000292" AFTER 06760 ns,
x"00000000" AFTER 06780 ns,
x"0000028E" AFTER 06800 ns,
x"00000000" AFTER 06820 ns,
x"0000028A" AFTER 06840 ns,
x"00000000" AFTER 06860 ns,
x"00000286" AFTER 06880 ns,
x"00000000" AFTER 06900 ns,
x"00000282" AFTER 06920 ns,
x"00000000" AFTER 06940 ns,
x"0000027E" AFTER 06960 ns,
x"00000000" AFTER 06980 ns,
x"0000027A" AFTER 07000 ns,
x"00000000" AFTER 07020 ns,
x"00000276" AFTER 07040 ns,
x"00000000" AFTER 07060 ns,
x"00000272" AFTER 07080 ns,
x"00000000" AFTER 07100 ns,
x"0000026E" AFTER 07120 ns,
x"00000000" AFTER 07140 ns,
x"0000026A" AFTER 07160 ns,
x"00000000" AFTER 07180 ns,
x"00000266" AFTER 07200 ns,
x"00000000" AFTER 07220 ns,
x"00000262" AFTER 07240 ns,
x"00000000" AFTER 07260 ns,
x"0000025E" AFTER 07280 ns,
x"00000000" AFTER 07300 ns,
x"0000025A" AFTER 07320 ns,
x"00000000" AFTER 07340 ns,
x"00000256" AFTER 07360 ns,
x"00000000" AFTER 07380 ns,
x"00000252" AFTER 07400 ns,
x"00000000" AFTER 07420 ns,
x"0000024E" AFTER 07440 ns,
x"00000000" AFTER 07460 ns,
x"0000024A" AFTER 07480 ns,
x"00000000" AFTER 07500 ns,
x"00000246" AFTER 07520 ns,
x"00000000" AFTER 07540 ns,
x"00000242" AFTER 07560 ns,
x"00000000" AFTER 07580 ns,
x"0000023E" AFTER 07600 ns,
x"00000000" AFTER 07620 ns,
x"0000023A" AFTER 07640 ns,
x"00000000" AFTER 07660 ns,
x"00000236" AFTER 07680 ns,
x"00000000" AFTER 07700 ns,
x"00000232" AFTER 07720 ns,
x"00000000" AFTER 07740 ns,
x"0000022E" AFTER 07760 ns,
x"00000000" AFTER 07780 ns,
x"0000022A" AFTER 07800 ns,
x"00000000" AFTER 07820 ns,
x"00000226" AFTER 07840 ns,
x"00000000" AFTER 07860 ns,
x"00000222" AFTER 07880 ns,
x"00000000" AFTER 07900 ns,
x"0000021E" AFTER 07920 ns,
x"00000000" AFTER 07940 ns,
x"0000021A" AFTER 07960 ns,
x"00000000" AFTER 07980 ns,
x"00000216" AFTER 08000 ns,
x"00000000" AFTER 08020 ns,
x"00000212" AFTER 08040 ns,
x"00000000" AFTER 08060 ns,
x"0000020E" AFTER 08080 ns,
x"00000000" AFTER 08100 ns,
x"0000020A" AFTER 08120 ns,
x"00000000" AFTER 08140 ns,
x"00000206" AFTER 08160 ns,
x"00000000" AFTER 08180 ns,
x"00000202" AFTER 08200 ns,
x"00000000" AFTER 08220 ns,
x"000001FE" AFTER 08240 ns,
x"00000000" AFTER 08260 ns,
x"000001FA" AFTER 08280 ns,
x"00000000" AFTER 08300 ns,
x"000001F6" AFTER 08320 ns,
x"00000000" AFTER 08340 ns,
x"000001F2" AFTER 08360 ns,
x"00000000" AFTER 08380 ns,
x"000001EE" AFTER 08400 ns,
x"00000000" AFTER 08420 ns,
x"000001EA" AFTER 08440 ns,
x"00000000" AFTER 08460 ns,
x"000001E6" AFTER 08480 ns,
x"00000000" AFTER 08500 ns,
x"000001E2" AFTER 08520 ns,
x"00000000" AFTER 08540 ns,
x"000001DE" AFTER 08560 ns,
x"00000000" AFTER 08580 ns,
x"000001DA" AFTER 08600 ns,
x"00000000" AFTER 08620 ns,
x"000001D6" AFTER 08640 ns,
x"00000000" AFTER 08660 ns,
x"000001D2" AFTER 08680 ns,
x"00000000" AFTER 08700 ns,
x"000001CE" AFTER 08720 ns,
x"00000000" AFTER 08740 ns,
x"000001CA" AFTER 08760 ns,
x"00000000" AFTER 08780 ns,
x"000001C6" AFTER 08800 ns,
x"00000000" AFTER 08820 ns,
x"000001C2" AFTER 08840 ns,
x"00000000" AFTER 08860 ns,
x"000001BE" AFTER 08880 ns,
x"00000000" AFTER 08900 ns,
x"000001BA" AFTER 08920 ns,
x"00000000" AFTER 08940 ns,
x"000001B6" AFTER 08960 ns,
x"00000000" AFTER 08980 ns,
x"000001B2" AFTER 09000 ns,
x"00000000" AFTER 09020 ns,
x"000001AE" AFTER 09040 ns,
x"00000000" AFTER 09060 ns,
x"000001AA" AFTER 09080 ns,
x"00000000" AFTER 09100 ns,
x"000001A6" AFTER 09120 ns,
x"00000000" AFTER 09140 ns,
x"000001A2" AFTER 09160 ns,
x"00000000" AFTER 09180 ns,
x"0000019E" AFTER 09200 ns,
x"00000000" AFTER 09220 ns,
x"0000019A" AFTER 09240 ns,
x"00000000" AFTER 09260 ns,
x"00000196" AFTER 09280 ns,
x"00000000" AFTER 09300 ns,
x"00000192" AFTER 09320 ns,
x"00000000" AFTER 09340 ns,
x"0000018E" AFTER 09360 ns,
x"00000000" AFTER 09380 ns,
x"0000018A" AFTER 09400 ns,
x"00000000" AFTER 09420 ns,
x"00000186" AFTER 09440 ns,
x"00000000" AFTER 09460 ns,
x"00000182" AFTER 09480 ns,
x"00000000" AFTER 09500 ns,
x"0000017E" AFTER 09520 ns,
x"00000000" AFTER 09540 ns,
x"0000017A" AFTER 09560 ns,
x"00000000" AFTER 09580 ns,
x"00000176" AFTER 09600 ns,
x"00000000" AFTER 09620 ns,
x"00000172" AFTER 09640 ns,
x"00000000" AFTER 09660 ns,
x"0000016E" AFTER 09680 ns,
x"00000000" AFTER 09700 ns,
x"0000016A" AFTER 09720 ns,
x"00000000" AFTER 09740 ns,
x"00000166" AFTER 09760 ns,
x"00000000" AFTER 09780 ns,
x"00000162" AFTER 09800 ns,
x"00000000" AFTER 09820 ns,
x"0000015E" AFTER 09840 ns,
x"00000000" AFTER 09860 ns,
x"0000015A" AFTER 09880 ns,
x"00000000" AFTER 09900 ns,
x"00000156" AFTER 09920 ns,
x"00000000" AFTER 09940 ns,
x"00000152" AFTER 09960 ns,
x"00000000" AFTER 09980 ns,
x"0000014E" AFTER 10000 ns,
x"00000000" AFTER 10020 ns,
x"0000014A" AFTER 10040 ns,
x"00000000" AFTER 10060 ns,
x"00000146" AFTER 10080 ns,
x"00000000" AFTER 10100 ns,
x"00000142" AFTER 10120 ns,
x"00000000" AFTER 10140 ns,
x"0000013E" AFTER 10160 ns,
x"00000000" AFTER 10180 ns,
x"0000013A" AFTER 10200 ns,
x"00000000" AFTER 10220 ns,
x"00000136" AFTER 10240 ns,
x"00000000" AFTER 10260 ns,
x"00000132" AFTER 10280 ns,
x"00000000" AFTER 10300 ns,
x"0000012E" AFTER 10320 ns,
x"00000000" AFTER 10340 ns,
x"0000012A" AFTER 10360 ns,
x"00000000" AFTER 10380 ns,
x"00000126" AFTER 10400 ns,
x"00000000" AFTER 10420 ns,
x"00000122" AFTER 10440 ns,
x"00000000" AFTER 10460 ns,
x"0000011E" AFTER 10480 ns,
x"00000000" AFTER 10500 ns,
x"0000011A" AFTER 10520 ns,
x"00000000" AFTER 10540 ns,
x"00000116" AFTER 10560 ns,
x"00000000" AFTER 10580 ns,
x"00000112" AFTER 10600 ns,
x"00000000" AFTER 10620 ns,
x"0000010E" AFTER 10640 ns,
x"00000000" AFTER 10660 ns,
x"0000010A" AFTER 10680 ns,
x"00000000" AFTER 10700 ns,
x"00000106" AFTER 10720 ns,
x"00000000" AFTER 10740 ns,
x"00000102" AFTER 10760 ns,
x"00000000" AFTER 10780 ns,
x"000000FE" AFTER 10800 ns,
x"00000000" AFTER 10820 ns,
x"000000FA" AFTER 10840 ns,
x"00000000" AFTER 10860 ns,
x"000000F6" AFTER 10880 ns,
x"00000000" AFTER 10900 ns,
x"000000F2" AFTER 10920 ns,
x"00000000" AFTER 10940 ns,
x"000000EE" AFTER 10960 ns,
x"00000000" AFTER 10980 ns,
x"000000EA" AFTER 11000 ns,
x"00000000" AFTER 11020 ns,
x"000000E6" AFTER 11040 ns,
x"00000000" AFTER 11060 ns,
x"000000E2" AFTER 11080 ns,
x"00000000" AFTER 11100 ns,
x"000000DE" AFTER 11120 ns,
x"00000000" AFTER 11140 ns,
x"000000DA" AFTER 11160 ns,
x"00000000" AFTER 11180 ns,
x"000000D6" AFTER 11200 ns,
x"00000000" AFTER 11220 ns,
x"000000D2" AFTER 11240 ns,
x"00000000" AFTER 11260 ns,
x"000000CE" AFTER 11280 ns,
x"00000000" AFTER 11300 ns,
x"000000CA" AFTER 11320 ns,
x"00000000" AFTER 11340 ns,
x"000000C6" AFTER 11360 ns,
x"00000000" AFTER 11380 ns,
x"000000C2" AFTER 11400 ns,
x"00000000" AFTER 11420 ns,
x"000000BE" AFTER 11440 ns,
x"00000000" AFTER 11460 ns,
x"000000BA" AFTER 11480 ns,
x"00000000" AFTER 11500 ns,
x"000000B6" AFTER 11520 ns,
x"00000000" AFTER 11540 ns,
x"000000B2" AFTER 11560 ns,
x"00000000" AFTER 11580 ns,
x"000000AE" AFTER 11600 ns,
x"00000000" AFTER 11620 ns,
x"000000AA" AFTER 11640 ns,
x"00000000" AFTER 11660 ns,
x"000000A6" AFTER 11680 ns,
x"00000000" AFTER 11700 ns,
x"000000A2" AFTER 11720 ns,
x"00000000" AFTER 11740 ns,
x"0000009E" AFTER 11760 ns,
x"00000000" AFTER 11780 ns,
x"0000009A" AFTER 11800 ns,
x"00000000" AFTER 11820 ns,
x"00000096" AFTER 11840 ns,
x"00000000" AFTER 11860 ns,
x"00000092" AFTER 11880 ns,
x"00000000" AFTER 11900 ns,
x"0000008E" AFTER 11920 ns,
x"00000000" AFTER 11940 ns,
x"0000008A" AFTER 11960 ns,
x"00000000" AFTER 11980 ns,
x"00000086" AFTER 12000 ns,
x"00000000" AFTER 12020 ns,
x"00000082" AFTER 12040 ns,
x"00000000" AFTER 12060 ns,
x"0000007E" AFTER 12080 ns,
x"00000000" AFTER 12100 ns,
x"0000007A" AFTER 12120 ns,
x"00000000" AFTER 12140 ns,
x"00000076" AFTER 12160 ns,
x"00000000" AFTER 12180 ns,
x"00000072" AFTER 12200 ns,
x"00000000" AFTER 12220 ns,
x"0000006E" AFTER 12240 ns,
x"00000000" AFTER 12260 ns,
x"0000006A" AFTER 12280 ns,
x"00000000" AFTER 12300 ns,
x"00000066" AFTER 12320 ns,
x"00000000" AFTER 12340 ns,
x"00000062" AFTER 12360 ns,
x"00000000" AFTER 12380 ns,
x"0000005E" AFTER 12400 ns,
x"00000000" AFTER 12420 ns,
x"0000005A" AFTER 12440 ns,
x"00000000" AFTER 12460 ns,
x"00000056" AFTER 12480 ns,
x"00000000" AFTER 12500 ns,
x"00000052" AFTER 12520 ns,
x"00000000" AFTER 12540 ns,
x"0000004E" AFTER 12560 ns,
x"00000000" AFTER 12580 ns,
x"0000004A" AFTER 12600 ns,
x"00000000" AFTER 12620 ns,
x"00000046" AFTER 12640 ns,
x"00000000" AFTER 12660 ns,
x"00000042" AFTER 12680 ns,
x"00000000" AFTER 12700 ns,
x"0000003E" AFTER 12720 ns,
x"00000000" AFTER 12740 ns,
x"0000003A" AFTER 12760 ns,
x"00000000" AFTER 12780 ns,
x"00000036" AFTER 12800 ns,
x"00000000" AFTER 12820 ns,
x"00000032" AFTER 12840 ns,
x"00000000" AFTER 12860 ns,
x"0000002E" AFTER 12880 ns,
x"00000000" AFTER 12900 ns,
x"0000002A" AFTER 12920 ns,
x"00000000" AFTER 12940 ns,
x"00000026" AFTER 12960 ns,
x"00000000" AFTER 12980 ns,
x"00000022" AFTER 13000 ns,
x"00000000" AFTER 13020 ns,
x"0000001E" AFTER 13040 ns,
x"00000000" AFTER 13060 ns,
x"0000001A" AFTER 13080 ns,
x"00000000" AFTER 13100 ns,
x"00000016" AFTER 13120 ns,
x"00000000" AFTER 13140 ns,
x"00000012" AFTER 13160 ns,
x"00000000" AFTER 13180 ns,
x"0000000E" AFTER 13200 ns,
x"00000000" AFTER 13220 ns,
x"0000000A" AFTER 13240 ns,
x"00000000" AFTER 13260 ns,
x"00000006" AFTER 13280 ns,
x"00000000" AFTER 13300 ns,
x"00000002" AFTER 13320 ns,
x"00000000" AFTER 13340 ns,
x"EE6B27FA" AFTER 13360 ns,
x"00000000" AFTER 13380 ns,
x"EE6B27F6" AFTER 13400 ns,
x"00000000" AFTER 13420 ns,
x"EE6B27F2" AFTER 13440 ns,
x"00000000" AFTER 13460 ns,
x"EE6B27EE" AFTER 13480 ns,
x"00000000" AFTER 13500 ns,
x"EE6B27EA" AFTER 13520 ns,
x"00000000" AFTER 13540 ns,
x"EE6B27E6" AFTER 13560 ns,
x"00000000" AFTER 13580 ns,
x"EE6B27E2" AFTER 13600 ns,
x"00000000" AFTER 13620 ns,
x"EE6B27DE" AFTER 13640 ns,
x"00000000" AFTER 13660 ns,
x"EE6B27DA" AFTER 13680 ns,
x"00000000" AFTER 13700 ns,
x"EE6B27D6" AFTER 13720 ns,
x"00000000" AFTER 13740 ns,
x"EE6B27D2" AFTER 13760 ns,
x"00000000" AFTER 13780 ns,
x"EE6B27CE" AFTER 13800 ns,
x"00000000" AFTER 13820 ns,
x"EE6B27CA" AFTER 13840 ns,
x"00000000" AFTER 13860 ns,
x"EE6B27C6" AFTER 13880 ns,
x"00000000" AFTER 13900 ns,
x"EE6B27C2" AFTER 13920 ns,
x"00000000" AFTER 13940 ns,
x"EE6B27BE" AFTER 13960 ns,
x"00000000" AFTER 13980 ns,
x"EE6B27BA" AFTER 14000 ns,
x"00000000" AFTER 14020 ns,
x"EE6B27B6" AFTER 14040 ns,
x"00000000" AFTER 14060 ns,
x"EE6B27B2" AFTER 14080 ns,
x"00000000" AFTER 14100 ns,
x"EE6B27AE" AFTER 14120 ns,
x"00000000" AFTER 14140 ns,
x"EE6B27AA" AFTER 14160 ns,
x"00000000" AFTER 14180 ns,
x"EE6B27A6" AFTER 14200 ns,
x"00000000" AFTER 14220 ns,
x"EE6B27A2" AFTER 14240 ns,
x"00000000" AFTER 14260 ns,
x"EE6B279E" AFTER 14280 ns,
x"00000000" AFTER 14300 ns,
x"EE6B279A" AFTER 14320 ns,
x"00000000" AFTER 14340 ns,
x"EE6B2796" AFTER 14360 ns,
x"00000000" AFTER 14380 ns,
x"EE6B2792" AFTER 14400 ns,
x"00000000" AFTER 14420 ns,
x"EE6B278E" AFTER 14440 ns,
x"00000000" AFTER 14460 ns,
x"EE6B278A" AFTER 14480 ns,
x"00000000" AFTER 14500 ns,
x"EE6B2786" AFTER 14520 ns,
x"00000000" AFTER 14540 ns,
x"EE6B2782" AFTER 14560 ns,
x"00000000" AFTER 14580 ns,
x"EE6B277E" AFTER 14600 ns,
x"00000000" AFTER 14620 ns,
x"EE6B277A" AFTER 14640 ns,
x"00000000" AFTER 14660 ns,
x"EE6B2776" AFTER 14680 ns,
x"00000000" AFTER 14700 ns,
x"EE6B2772" AFTER 14720 ns,
x"00000000" AFTER 14740 ns,
x"EE6B276E" AFTER 14760 ns,
x"00000000" AFTER 14780 ns,
x"EE6B276A" AFTER 14800 ns,
x"00000000" AFTER 14820 ns,
x"EE6B2766" AFTER 14840 ns,
x"00000000" AFTER 14860 ns,
x"EE6B2762" AFTER 14880 ns,
x"00000000" AFTER 14900 ns,
x"EE6B275E" AFTER 14920 ns,
x"00000000" AFTER 14940 ns,
x"EE6B275A" AFTER 14960 ns,
x"00000000" AFTER 14980 ns,
x"EE6B2756" AFTER 15000 ns,
x"00000000" AFTER 15020 ns,
x"EE6B2752" AFTER 15040 ns,
x"00000000" AFTER 15060 ns,
x"EE6B274E" AFTER 15080 ns,
x"00000000" AFTER 15100 ns,
x"EE6B274A" AFTER 15120 ns,
x"00000000" AFTER 15140 ns,
x"EE6B2746" AFTER 15160 ns,
x"00000000" AFTER 15180 ns,
x"EE6B2742" AFTER 15200 ns,
x"00000000" AFTER 15220 ns,
x"EE6B273E" AFTER 15240 ns,
x"00000000" AFTER 15260 ns,
x"EE6B273A" AFTER 15280 ns,
x"00000000" AFTER 15300 ns,
x"EE6B2736" AFTER 15320 ns,
x"00000000" AFTER 15340 ns,
x"EE6B2732" AFTER 15360 ns,
x"00000000" AFTER 15380 ns,
x"EE6B272E" AFTER 15400 ns,
x"00000000" AFTER 15420 ns,
x"EE6B272A" AFTER 15440 ns,
x"00000000" AFTER 15460 ns,
x"EE6B2726" AFTER 15480 ns,
x"00000000" AFTER 15500 ns,
x"EE6B2722" AFTER 15520 ns,
x"00000000" AFTER 15540 ns,
x"EE6B271E" AFTER 15560 ns,
x"00000000" AFTER 15580 ns,
x"EE6B271A" AFTER 15600 ns,
x"00000000" AFTER 15620 ns,
x"EE6B2716" AFTER 15640 ns,
x"00000000" AFTER 15660 ns,
x"EE6B2712" AFTER 15680 ns,
x"00000000" AFTER 15700 ns,
x"EE6B270E" AFTER 15720 ns,
x"00000000" AFTER 15740 ns,
x"EE6B270A" AFTER 15760 ns,
x"00000000" AFTER 15780 ns,
x"EE6B2706" AFTER 15800 ns,
x"00000000" AFTER 15820 ns,
x"EE6B2702" AFTER 15840 ns,
x"00000000" AFTER 15860 ns,
x"EE6B26FE" AFTER 15880 ns,
x"00000000" AFTER 15900 ns,
x"EE6B26FA" AFTER 15920 ns,
x"00000000" AFTER 15940 ns,
x"EE6B26F6" AFTER 15960 ns,
x"00000000" AFTER 15980 ns,
x"EE6B26F2" AFTER 16000 ns,
x"00000000" AFTER 16020 ns,
x"EE6B26EE" AFTER 16040 ns,
x"00000000" AFTER 16060 ns,
x"EE6B26EA" AFTER 16080 ns,
x"00000000" AFTER 16100 ns,
x"EE6B26E6" AFTER 16120 ns,
x"00000000" AFTER 16140 ns,
x"EE6B26E2" AFTER 16160 ns,
x"00000000" AFTER 16180 ns,
x"EE6B26DE" AFTER 16200 ns,
x"00000000" AFTER 16220 ns,
x"EE6B26DA" AFTER 16240 ns,
x"00000000" AFTER 16260 ns,
x"EE6B26D6" AFTER 16280 ns,
x"00000000" AFTER 16300 ns,
x"EE6B26D2" AFTER 16320 ns,
x"00000000" AFTER 16340 ns,
x"EE6B26CE" AFTER 16360 ns,
x"00000000" AFTER 16380 ns,
x"EE6B26CA" AFTER 16400 ns,
x"00000000" AFTER 16420 ns,
x"EE6B26C6" AFTER 16440 ns,
x"00000000" AFTER 16460 ns,
x"EE6B26C2" AFTER 16480 ns,
x"00000000" AFTER 16500 ns,
x"EE6B26BE" AFTER 16520 ns,
x"00000000" AFTER 16540 ns,
x"EE6B26BA" AFTER 16560 ns,
x"00000000" AFTER 16580 ns,
x"EE6B26B6" AFTER 16600 ns,
x"00000000" AFTER 16620 ns,
x"EE6B26B2" AFTER 16640 ns,
x"00000000" AFTER 16660 ns,
x"EE6B26AE" AFTER 16680 ns,
x"00000000" AFTER 16700 ns,
x"EE6B26AA" AFTER 16720 ns,
x"00000000" AFTER 16740 ns,
x"EE6B26A6" AFTER 16760 ns,
x"00000000" AFTER 16780 ns,
x"EE6B26A2" AFTER 16800 ns,
x"00000000" AFTER 16820 ns,
x"EE6B269E" AFTER 16840 ns,
x"00000000" AFTER 16860 ns,
x"EE6B269A" AFTER 16880 ns,
x"00000000" AFTER 16900 ns,
x"EE6B2696" AFTER 16920 ns,
x"00000000" AFTER 16940 ns,
x"EE6B2692" AFTER 16960 ns,
x"00000000" AFTER 16980 ns,
x"EE6B268E" AFTER 17000 ns,
x"00000000" AFTER 17020 ns,
x"EE6B268A" AFTER 17040 ns,
x"00000000" AFTER 17060 ns,
x"EE6B2686" AFTER 17080 ns,
x"00000000" AFTER 17100 ns,
x"EE6B2682" AFTER 17120 ns,
x"00000000" AFTER 17140 ns,
x"EE6B267E" AFTER 17160 ns,
x"00000000" AFTER 17180 ns,
x"EE6B267A" AFTER 17200 ns,
x"00000000" AFTER 17220 ns,
x"EE6B2676" AFTER 17240 ns,
x"00000000" AFTER 17260 ns,
x"EE6B2672" AFTER 17280 ns,
x"00000000" AFTER 17300 ns,
x"EE6B266E" AFTER 17320 ns,
x"00000000" AFTER 17340 ns,
x"EE6B266A" AFTER 17360 ns,
x"00000000" AFTER 17380 ns,
x"EE6B2666" AFTER 17400 ns,
x"00000000" AFTER 17420 ns,
x"EE6B2662" AFTER 17440 ns,
x"00000000" AFTER 17460 ns,
x"EE6B265E" AFTER 17480 ns,
x"00000000" AFTER 17500 ns,
x"EE6B265A" AFTER 17520 ns,
x"00000000" AFTER 17540 ns,
x"EE6B2656" AFTER 17560 ns,
x"00000000" AFTER 17580 ns,
x"EE6B2652" AFTER 17600 ns,
x"00000000" AFTER 17620 ns,
x"EE6B264E" AFTER 17640 ns,
x"00000000" AFTER 17660 ns,
x"EE6B264A" AFTER 17680 ns,
x"00000000" AFTER 17700 ns,
x"EE6B2646" AFTER 17720 ns,
x"00000000" AFTER 17740 ns,
x"EE6B2642" AFTER 17760 ns,
x"00000000" AFTER 17780 ns,
x"EE6B263E" AFTER 17800 ns,
x"00000000" AFTER 17820 ns,
x"EE6B263A" AFTER 17840 ns,
x"00000000" AFTER 17860 ns,
x"EE6B2636" AFTER 17880 ns,
x"00000000" AFTER 17900 ns,
x"EE6B2632" AFTER 17920 ns,
x"00000000" AFTER 17940 ns,
x"EE6B262E" AFTER 17960 ns,
x"00000000" AFTER 17980 ns,
x"EE6B262A" AFTER 18000 ns,
x"00000000" AFTER 18020 ns,
x"EE6B2626" AFTER 18040 ns,
x"00000000" AFTER 18060 ns,
x"EE6B2622" AFTER 18080 ns,
x"00000000" AFTER 18100 ns,
x"EE6B261E" AFTER 18120 ns,
x"00000000" AFTER 18140 ns,
x"EE6B261A" AFTER 18160 ns,
x"00000000" AFTER 18180 ns,
x"EE6B2616" AFTER 18200 ns,
x"00000000" AFTER 18220 ns,
x"EE6B2612" AFTER 18240 ns,
x"00000000" AFTER 18260 ns,
x"EE6B260E" AFTER 18280 ns,
x"00000000" AFTER 18300 ns,
x"EE6B260A" AFTER 18320 ns,
x"00000000" AFTER 18340 ns,
x"EE6B2606" AFTER 18360 ns,
x"00000000" AFTER 18380 ns,
x"EE6B2602" AFTER 18400 ns,
x"00000000" AFTER 18420 ns,
x"EE6B25FE" AFTER 18440 ns,
x"00000000" AFTER 18460 ns,
x"EE6B25FA" AFTER 18480 ns,
x"00000000" AFTER 18500 ns,
x"EE6B25F6" AFTER 18520 ns,
x"00000000" AFTER 18540 ns,
x"EE6B25F2" AFTER 18560 ns,
x"00000000" AFTER 18580 ns,
x"EE6B25EE" AFTER 18600 ns,
x"00000000" AFTER 18620 ns,
x"EE6B25EA" AFTER 18640 ns,
x"00000000" AFTER 18660 ns,
x"EE6B25E6" AFTER 18680 ns,
x"00000000" AFTER 18700 ns,
x"EE6B25E2" AFTER 18720 ns,
x"00000000" AFTER 18740 ns,
x"EE6B25DE" AFTER 18760 ns,
x"00000000" AFTER 18780 ns,
x"EE6B25DA" AFTER 18800 ns,
x"00000000" AFTER 18820 ns,
x"EE6B25D6" AFTER 18840 ns,
x"00000000" AFTER 18860 ns,
x"EE6B25D2" AFTER 18880 ns,
x"00000000" AFTER 18900 ns,
x"EE6B25CE" AFTER 18920 ns,
x"00000000" AFTER 18940 ns,
x"EE6B25CA" AFTER 18960 ns,
x"00000000" AFTER 18980 ns,
x"EE6B25C6" AFTER 19000 ns,
x"00000000" AFTER 19020 ns,
x"EE6B25C2" AFTER 19040 ns,
x"00000000" AFTER 19060 ns,
x"EE6B25BE" AFTER 19080 ns,
x"00000000" AFTER 19100 ns,
x"EE6B25BA" AFTER 19120 ns,
x"00000000" AFTER 19140 ns,
x"EE6B25B6" AFTER 19160 ns,
x"00000000" AFTER 19180 ns,
x"EE6B25B2" AFTER 19200 ns,
x"00000000" AFTER 19220 ns,
x"EE6B25AE" AFTER 19240 ns,
x"00000000" AFTER 19260 ns,
x"EE6B25AA" AFTER 19280 ns,
x"00000000" AFTER 19300 ns,
x"EE6B25A6" AFTER 19320 ns,
x"00000000" AFTER 19340 ns,
x"EE6B25A2" AFTER 19360 ns,
x"00000000" AFTER 19380 ns,
x"EE6B259E" AFTER 19400 ns,
x"00000000" AFTER 19420 ns,
x"EE6B259A" AFTER 19440 ns,
x"00000000" AFTER 19460 ns,
x"EE6B2596" AFTER 19480 ns,
x"00000000" AFTER 19500 ns,
x"EE6B2592" AFTER 19520 ns,
x"00000000" AFTER 19540 ns,
x"EE6B258E" AFTER 19560 ns,
x"00000000" AFTER 19580 ns,
x"EE6B258A" AFTER 19600 ns,
x"00000000" AFTER 19620 ns,
x"EE6B2586" AFTER 19640 ns,
x"00000000" AFTER 19660 ns,
x"EE6B2582" AFTER 19680 ns,
x"00000000" AFTER 19700 ns,
x"EE6B257E" AFTER 19720 ns,
x"00000000" AFTER 19740 ns,
x"EE6B257A" AFTER 19760 ns,
x"00000000" AFTER 19780 ns,
x"EE6B2576" AFTER 19800 ns,
x"00000000" AFTER 19820 ns,
x"EE6B2572" AFTER 19840 ns,
x"00000000" AFTER 19860 ns,
x"EE6B256E" AFTER 19880 ns,
x"00000000" AFTER 19900 ns,
x"EE6B256A" AFTER 19920 ns,
x"00000000" AFTER 19940 ns,
x"EE6B256E" AFTER 19960 ns,
x"00000000" AFTER 19980 ns,
x"EE6B2572" AFTER 20000 ns,
x"00000000" AFTER 20020 ns,
x"EE6B2576" AFTER 20040 ns,
x"00000000" AFTER 20060 ns,
x"EE6B257A" AFTER 20080 ns,
x"00000000" AFTER 20100 ns,
x"EE6B257E" AFTER 20120 ns,
x"00000000" AFTER 20140 ns,
x"EE6B2582" AFTER 20160 ns,
x"00000000" AFTER 20180 ns,
x"EE6B2586" AFTER 20200 ns,
x"00000000" AFTER 20220 ns,
x"EE6B258A" AFTER 20240 ns,
x"00000000" AFTER 20260 ns,
x"EE6B258E" AFTER 20280 ns,
x"00000000" AFTER 20300 ns,
x"EE6B2592" AFTER 20320 ns,
x"00000000" AFTER 20340 ns,
x"EE6B2596" AFTER 20360 ns,
x"00000000" AFTER 20380 ns,
x"EE6B259A" AFTER 20400 ns,
x"00000000" AFTER 20420 ns,
x"EE6B259E" AFTER 20440 ns,
x"00000000" AFTER 20460 ns,
x"EE6B25A2" AFTER 20480 ns,
x"00000000" AFTER 20500 ns,
x"EE6B25A6" AFTER 20520 ns,
x"00000000" AFTER 20540 ns,
x"EE6B25AA" AFTER 20560 ns,
x"00000000" AFTER 20580 ns,
x"EE6B25AE" AFTER 20600 ns,
x"00000000" AFTER 20620 ns,
x"EE6B25B2" AFTER 20640 ns,
x"00000000" AFTER 20660 ns,
x"EE6B25B6" AFTER 20680 ns,
x"00000000" AFTER 20700 ns,
x"EE6B25BA" AFTER 20720 ns,
x"00000000" AFTER 20740 ns,
x"EE6B25BE" AFTER 20760 ns,
x"00000000" AFTER 20780 ns,
x"EE6B25C2" AFTER 20800 ns,
x"00000000" AFTER 20820 ns,
x"EE6B25C6" AFTER 20840 ns,
x"00000000" AFTER 20860 ns,
x"EE6B25CA" AFTER 20880 ns,
x"00000000" AFTER 20900 ns,
x"EE6B25CE" AFTER 20920 ns,
x"00000000" AFTER 20940 ns,
x"EE6B25D2" AFTER 20960 ns,
x"00000000" AFTER 20980 ns,
x"EE6B25D6" AFTER 21000 ns,
x"00000000" AFTER 21020 ns,
x"EE6B25DA" AFTER 21040 ns,
x"00000000" AFTER 21060 ns,
x"EE6B25DE" AFTER 21080 ns,
x"00000000" AFTER 21100 ns,
x"EE6B25E2" AFTER 21120 ns,
x"00000000" AFTER 21140 ns,
x"EE6B25E6" AFTER 21160 ns,
x"00000000" AFTER 21180 ns,
x"EE6B25EA" AFTER 21200 ns,
x"00000000" AFTER 21220 ns,
x"EE6B25EE" AFTER 21240 ns,
x"00000000" AFTER 21260 ns,
x"EE6B25F2" AFTER 21280 ns,
x"00000000" AFTER 21300 ns,
x"EE6B25F6" AFTER 21320 ns,
x"00000000" AFTER 21340 ns,
x"EE6B25FA" AFTER 21360 ns,
x"00000000" AFTER 21380 ns,
x"EE6B25FE" AFTER 21400 ns,
x"00000000" AFTER 21420 ns,
x"EE6B2602" AFTER 21440 ns,
x"00000000" AFTER 21460 ns,
x"EE6B2606" AFTER 21480 ns,
x"00000000" AFTER 21500 ns,
x"EE6B260A" AFTER 21520 ns,
x"00000000" AFTER 21540 ns,
x"EE6B260E" AFTER 21560 ns,
x"00000000" AFTER 21580 ns,
x"EE6B2612" AFTER 21600 ns,
x"00000000" AFTER 21620 ns,
x"EE6B2616" AFTER 21640 ns,
x"00000000" AFTER 21660 ns,
x"EE6B261A" AFTER 21680 ns,
x"00000000" AFTER 21700 ns,
x"EE6B261E" AFTER 21720 ns,
x"00000000" AFTER 21740 ns,
x"EE6B2622" AFTER 21760 ns,
x"00000000" AFTER 21780 ns,
x"EE6B2626" AFTER 21800 ns,
x"00000000" AFTER 21820 ns,
x"EE6B262A" AFTER 21840 ns,
x"00000000" AFTER 21860 ns,
x"EE6B262E" AFTER 21880 ns,
x"00000000" AFTER 21900 ns,
x"EE6B2632" AFTER 21920 ns,
x"00000000" AFTER 21940 ns,
x"EE6B2636" AFTER 21960 ns,
x"00000000" AFTER 21980 ns,
x"EE6B263A" AFTER 22000 ns,
x"00000000" AFTER 22020 ns,
x"EE6B263E" AFTER 22040 ns,
x"00000000" AFTER 22060 ns,
x"EE6B2642" AFTER 22080 ns,
x"00000000" AFTER 22100 ns,
x"EE6B2646" AFTER 22120 ns,
x"00000000" AFTER 22140 ns,
x"EE6B264A" AFTER 22160 ns,
x"00000000" AFTER 22180 ns,
x"EE6B264E" AFTER 22200 ns,
x"00000000" AFTER 22220 ns,
x"EE6B2652" AFTER 22240 ns,
x"00000000" AFTER 22260 ns,
x"EE6B2656" AFTER 22280 ns,
x"00000000" AFTER 22300 ns,
x"EE6B265A" AFTER 22320 ns,
x"00000000" AFTER 22340 ns,
x"EE6B265E" AFTER 22360 ns,
x"00000000" AFTER 22380 ns,
x"EE6B2662" AFTER 22400 ns,
x"00000000" AFTER 22420 ns,
x"EE6B2666" AFTER 22440 ns,
x"00000000" AFTER 22460 ns,
x"EE6B266A" AFTER 22480 ns,
x"00000000" AFTER 22500 ns,
x"EE6B266E" AFTER 22520 ns,
x"00000000" AFTER 22540 ns,
x"EE6B2672" AFTER 22560 ns,
x"00000000" AFTER 22580 ns,
x"EE6B2676" AFTER 22600 ns,
x"00000000" AFTER 22620 ns,
x"EE6B267A" AFTER 22640 ns,
x"00000000" AFTER 22660 ns,
x"EE6B267E" AFTER 22680 ns,
x"00000000" AFTER 22700 ns,
x"EE6B2682" AFTER 22720 ns,
x"00000000" AFTER 22740 ns,
x"EE6B2686" AFTER 22760 ns,
x"00000000" AFTER 22780 ns,
x"EE6B268A" AFTER 22800 ns,
x"00000000" AFTER 22820 ns,
x"EE6B268E" AFTER 22840 ns,
x"00000000" AFTER 22860 ns,
x"EE6B2692" AFTER 22880 ns,
x"00000000" AFTER 22900 ns,
x"EE6B2696" AFTER 22920 ns,
x"00000000" AFTER 22940 ns,
x"EE6B269A" AFTER 22960 ns,
x"00000000" AFTER 22980 ns,
x"EE6B269E" AFTER 23000 ns,
x"00000000" AFTER 23020 ns,
x"EE6B26A2" AFTER 23040 ns,
x"00000000" AFTER 23060 ns,
x"EE6B26A6" AFTER 23080 ns,
x"00000000" AFTER 23100 ns,
x"EE6B26AA" AFTER 23120 ns,
x"00000000" AFTER 23140 ns,
x"EE6B26AE" AFTER 23160 ns,
x"00000000" AFTER 23180 ns,
x"EE6B26B2" AFTER 23200 ns,
x"00000000" AFTER 23220 ns,
x"EE6B26B6" AFTER 23240 ns,
x"00000000" AFTER 23260 ns,
x"EE6B26BA" AFTER 23280 ns,
x"00000000" AFTER 23300 ns,
x"EE6B26BE" AFTER 23320 ns,
x"00000000" AFTER 23340 ns,
x"EE6B26C2" AFTER 23360 ns,
x"00000000" AFTER 23380 ns,
x"EE6B26C6" AFTER 23400 ns,
x"00000000" AFTER 23420 ns,
x"EE6B26CA" AFTER 23440 ns,
x"00000000" AFTER 23460 ns,
x"EE6B26CE" AFTER 23480 ns,
x"00000000" AFTER 23500 ns,
x"EE6B26D2" AFTER 23520 ns,
x"00000000" AFTER 23540 ns,
x"EE6B26D6" AFTER 23560 ns,
x"00000000" AFTER 23580 ns,
x"EE6B26DA" AFTER 23600 ns,
x"00000000" AFTER 23620 ns,
x"EE6B26DE" AFTER 23640 ns,
x"00000000" AFTER 23660 ns,
x"EE6B26E2" AFTER 23680 ns,
x"00000000" AFTER 23700 ns,
x"EE6B26E6" AFTER 23720 ns,
x"00000000" AFTER 23740 ns,
x"EE6B26EA" AFTER 23760 ns,
x"00000000" AFTER 23780 ns,
x"EE6B26EE" AFTER 23800 ns,
x"00000000" AFTER 23820 ns,
x"EE6B26F2" AFTER 23840 ns,
x"00000000" AFTER 23860 ns,
x"EE6B26F6" AFTER 23880 ns,
x"00000000" AFTER 23900 ns,
x"EE6B26FA" AFTER 23920 ns,
x"00000000" AFTER 23940 ns,
x"EE6B26FE" AFTER 23960 ns,
x"00000000" AFTER 23980 ns,
x"EE6B2702" AFTER 24000 ns,
x"00000000" AFTER 24020 ns,
x"EE6B2706" AFTER 24040 ns,
x"00000000" AFTER 24060 ns,
x"EE6B270A" AFTER 24080 ns,
x"00000000" AFTER 24100 ns,
x"EE6B270E" AFTER 24120 ns,
x"00000000" AFTER 24140 ns,
x"EE6B2712" AFTER 24160 ns,
x"00000000" AFTER 24180 ns,
x"EE6B2716" AFTER 24200 ns,
x"00000000" AFTER 24220 ns,
x"EE6B271A" AFTER 24240 ns,
x"00000000" AFTER 24260 ns,
x"EE6B271E" AFTER 24280 ns,
x"00000000" AFTER 24300 ns,
x"EE6B2722" AFTER 24320 ns,
x"00000000" AFTER 24340 ns,
x"EE6B2726" AFTER 24360 ns,
x"00000000" AFTER 24380 ns,
x"EE6B272A" AFTER 24400 ns,
x"00000000" AFTER 24420 ns,
x"EE6B272E" AFTER 24440 ns,
x"00000000" AFTER 24460 ns,
x"EE6B2732" AFTER 24480 ns,
x"00000000" AFTER 24500 ns,
x"EE6B2736" AFTER 24520 ns,
x"00000000" AFTER 24540 ns,
x"EE6B273A" AFTER 24560 ns,
x"00000000" AFTER 24580 ns,
x"EE6B273E" AFTER 24600 ns,
x"00000000" AFTER 24620 ns,
x"EE6B2742" AFTER 24640 ns,
x"00000000" AFTER 24660 ns,
x"EE6B2746" AFTER 24680 ns,
x"00000000" AFTER 24700 ns,
x"EE6B274A" AFTER 24720 ns,
x"00000000" AFTER 24740 ns,
x"EE6B274E" AFTER 24760 ns,
x"00000000" AFTER 24780 ns,
x"EE6B2752" AFTER 24800 ns,
x"00000000" AFTER 24820 ns,
x"EE6B2756" AFTER 24840 ns,
x"00000000" AFTER 24860 ns,
x"EE6B275A" AFTER 24880 ns,
x"00000000" AFTER 24900 ns,
x"EE6B275E" AFTER 24920 ns,
x"00000000" AFTER 24940 ns,
x"EE6B2762" AFTER 24960 ns,
x"00000000" AFTER 24980 ns,
x"EE6B2766" AFTER 25000 ns,
x"00000000" AFTER 25020 ns,
x"EE6B276A" AFTER 25040 ns,
x"00000000" AFTER 25060 ns,
x"EE6B276E" AFTER 25080 ns,
x"00000000" AFTER 25100 ns,
x"EE6B2772" AFTER 25120 ns,
x"00000000" AFTER 25140 ns,
x"EE6B2776" AFTER 25160 ns,
x"00000000" AFTER 25180 ns,
x"EE6B277A" AFTER 25200 ns,
x"00000000" AFTER 25220 ns,
x"EE6B277E" AFTER 25240 ns,
x"00000000" AFTER 25260 ns,
x"EE6B2782" AFTER 25280 ns,
x"00000000" AFTER 25300 ns,
x"EE6B2786" AFTER 25320 ns,
x"00000000" AFTER 25340 ns,
x"EE6B278A" AFTER 25360 ns,
x"00000000" AFTER 25380 ns,
x"EE6B278E" AFTER 25400 ns,
x"00000000" AFTER 25420 ns,
x"EE6B2792" AFTER 25440 ns,
x"00000000" AFTER 25460 ns,
x"EE6B2796" AFTER 25480 ns,
x"00000000" AFTER 25500 ns,
x"EE6B279A" AFTER 25520 ns,
x"00000000" AFTER 25540 ns,
x"EE6B279E" AFTER 25560 ns,
x"00000000" AFTER 25580 ns,
x"EE6B27A2" AFTER 25600 ns,
x"00000000" AFTER 25620 ns,
x"EE6B27A6" AFTER 25640 ns,
x"00000000" AFTER 25660 ns,
x"EE6B27AA" AFTER 25680 ns,
x"00000000" AFTER 25700 ns,
x"EE6B27AE" AFTER 25720 ns,
x"00000000" AFTER 25740 ns,
x"EE6B27B2" AFTER 25760 ns,
x"00000000" AFTER 25780 ns,
x"EE6B27B6" AFTER 25800 ns,
x"00000000" AFTER 25820 ns,
x"EE6B27BA" AFTER 25840 ns,
x"00000000" AFTER 25860 ns,
x"EE6B27BE" AFTER 25880 ns,
x"00000000" AFTER 25900 ns,
x"EE6B27C2" AFTER 25920 ns,
x"00000000" AFTER 25940 ns,
x"EE6B27C6" AFTER 25960 ns,
x"00000000" AFTER 25980 ns,
x"EE6B27CA" AFTER 26000 ns,
x"00000000" AFTER 26020 ns,
x"EE6B27CE" AFTER 26040 ns,
x"00000000" AFTER 26060 ns,
x"EE6B27D2" AFTER 26080 ns,
x"00000000" AFTER 26100 ns,
x"EE6B27D6" AFTER 26120 ns,
x"00000000" AFTER 26140 ns,
x"EE6B27DA" AFTER 26160 ns,
x"00000000" AFTER 26180 ns,
x"EE6B27DE" AFTER 26200 ns,
x"00000000" AFTER 26220 ns,
x"EE6B27E2" AFTER 26240 ns,
x"00000000" AFTER 26260 ns,
x"EE6B27E6" AFTER 26280 ns,
x"00000000" AFTER 26300 ns,
x"EE6B27EA" AFTER 26320 ns,
x"00000000" AFTER 26340 ns,
x"EE6B27EE" AFTER 26360 ns,
x"00000000" AFTER 26380 ns,
x"EE6B27F2" AFTER 26400 ns,
x"00000000" AFTER 26420 ns,
x"EE6B27F6" AFTER 26440 ns,
x"00000000" AFTER 26460 ns,
x"EE6B27FA" AFTER 26480 ns,
x"00000000" AFTER 26500 ns,
x"EE6B27FE" AFTER 26520 ns,
x"00000000" AFTER 26540 ns,
x"EE6B2802" AFTER 26560 ns,
x"00000000" AFTER 26580 ns,
x"EE6B2806" AFTER 26600 ns,
x"00000000" AFTER 26620 ns,
x"EE6B280A" AFTER 26640 ns,
x"00000000" AFTER 26660 ns,
x"EE6B280E" AFTER 26680 ns,
x"00000000" AFTER 26700 ns,
x"EE6B2812" AFTER 26720 ns,
x"00000000" AFTER 26740 ns,
x"EE6B2816" AFTER 26760 ns,
x"00000000" AFTER 26780 ns,
x"EE6B281A" AFTER 26800 ns,
x"00000000" AFTER 26820 ns,
x"EE6B281E" AFTER 26840 ns,
x"00000000" AFTER 26860 ns,
x"EE6B2822" AFTER 26880 ns,
x"00000000" AFTER 26900 ns,
x"EE6B2826" AFTER 26920 ns,
x"00000000" AFTER 26940 ns,
x"EE6B282A" AFTER 26960 ns,
x"00000000" AFTER 26980 ns,
x"EE6B282E" AFTER 27000 ns,
x"00000000" AFTER 27020 ns,
x"EE6B2832" AFTER 27040 ns,
x"00000000" AFTER 27060 ns,
x"EE6B2836" AFTER 27080 ns,
x"00000000" AFTER 27100 ns,
x"EE6B283A" AFTER 27120 ns,
x"00000000" AFTER 27140 ns,
x"EE6B283E" AFTER 27160 ns,
x"00000000" AFTER 27180 ns,
x"EE6B2842" AFTER 27200 ns,
x"00000000" AFTER 27220 ns,
x"EE6B2846" AFTER 27240 ns,
x"00000000" AFTER 27260 ns,
x"EE6B284A" AFTER 27280 ns,
x"00000000" AFTER 27300 ns,
x"EE6B284E" AFTER 27320 ns,
x"00000000" AFTER 27340 ns,
x"EE6B2852" AFTER 27360 ns,
x"00000000" AFTER 27380 ns,
x"EE6B2856" AFTER 27400 ns,
x"00000000" AFTER 27420 ns,
x"EE6B285A" AFTER 27440 ns,
x"00000000" AFTER 27460 ns,
x"EE6B285E" AFTER 27480 ns,
x"00000000" AFTER 27500 ns,
x"EE6B2862" AFTER 27520 ns,
x"00000000" AFTER 27540 ns,
x"EE6B2866" AFTER 27560 ns,
x"00000000" AFTER 27580 ns,
x"EE6B286A" AFTER 27600 ns,
x"00000000" AFTER 27620 ns,
x"EE6B286E" AFTER 27640 ns,
x"00000000" AFTER 27660 ns,
x"EE6B2872" AFTER 27680 ns,
x"00000000" AFTER 27700 ns,
x"EE6B2876" AFTER 27720 ns,
x"00000000" AFTER 27740 ns,
x"EE6B287A" AFTER 27760 ns,
x"00000000" AFTER 27780 ns,
x"EE6B287E" AFTER 27800 ns,
x"00000000" AFTER 27820 ns,
x"EE6B2882" AFTER 27840 ns,
x"00000000" AFTER 27860 ns,
x"EE6B2886" AFTER 27880 ns,
x"00000000" AFTER 27900 ns,
x"EE6B288A" AFTER 27920 ns,
x"00000000" AFTER 27940 ns,
x"EE6B288E" AFTER 27960 ns,
x"00000000" AFTER 27980 ns,
x"EE6B2892" AFTER 28000 ns,
x"00000000" AFTER 28020 ns,
x"EE6B2896" AFTER 28040 ns,
x"00000000" AFTER 28060 ns,
x"EE6B289A" AFTER 28080 ns,
x"00000000" AFTER 28100 ns,
x"EE6B289E" AFTER 28120 ns,
x"00000000" AFTER 28140 ns,
x"EE6B28A2" AFTER 28160 ns,
x"00000000" AFTER 28180 ns,
x"EE6B28A6" AFTER 28200 ns,
x"00000000" AFTER 28220 ns,
x"EE6B28AA" AFTER 28240 ns,
x"00000000" AFTER 28260 ns,
x"EE6B28AE" AFTER 28280 ns,
x"00000000" AFTER 28300 ns,
x"EE6B28B2" AFTER 28320 ns,
x"00000000" AFTER 28340 ns,
x"EE6B28B6" AFTER 28360 ns,
x"00000000" AFTER 28380 ns,
x"EE6B28BA" AFTER 28400 ns,
x"00000000" AFTER 28420 ns,
x"EE6B28BE" AFTER 28440 ns,
x"00000000" AFTER 28460 ns,
x"EE6B28C2" AFTER 28480 ns,
x"00000000" AFTER 28500 ns,
x"EE6B28C6" AFTER 28520 ns,
x"00000000" AFTER 28540 ns,
x"EE6B28CA" AFTER 28560 ns,
x"00000000" AFTER 28580 ns,
x"EE6B28CE" AFTER 28600 ns,
x"00000000" AFTER 28620 ns,
x"EE6B28D2" AFTER 28640 ns,
x"00000000" AFTER 28660 ns,
x"EE6B28D6" AFTER 28680 ns,
x"00000000" AFTER 28700 ns,
x"EE6B28DA" AFTER 28720 ns,
x"00000000" AFTER 28740 ns,
x"EE6B28DE" AFTER 28760 ns,
x"00000000" AFTER 28780 ns,
x"EE6B28E2" AFTER 28800 ns,
x"00000000" AFTER 28820 ns,
x"EE6B28E6" AFTER 28840 ns,
x"00000000" AFTER 28860 ns,
x"EE6B28EA" AFTER 28880 ns,
x"00000000" AFTER 28900 ns,
x"EE6B28EE" AFTER 28920 ns,
x"00000000" AFTER 28940 ns,
x"EE6B28F2" AFTER 28960 ns,
x"00000000" AFTER 28980 ns,
x"EE6B28F6" AFTER 29000 ns,
x"00000000" AFTER 29020 ns,
x"EE6B28FA" AFTER 29040 ns,
x"00000000" AFTER 29060 ns,
x"EE6B28FE" AFTER 29080 ns,
x"00000000" AFTER 29100 ns,
x"EE6B2902" AFTER 29120 ns,
x"00000000" AFTER 29140 ns,
x"EE6B2906" AFTER 29160 ns,
x"00000000" AFTER 29180 ns,
x"EE6B290A" AFTER 29200 ns,
x"00000000" AFTER 29220 ns,
x"EE6B290E" AFTER 29240 ns,
x"00000000" AFTER 29260 ns,
x"EE6B2912" AFTER 29280 ns,
x"00000000" AFTER 29300 ns,
x"EE6B2916" AFTER 29320 ns,
x"00000000" AFTER 29340 ns,
x"EE6B291A" AFTER 29360 ns,
x"00000000" AFTER 29380 ns,
x"EE6B291E" AFTER 29400 ns,
x"00000000" AFTER 29420 ns,
x"EE6B2922" AFTER 29440 ns,
x"00000000" AFTER 29460 ns,
x"EE6B2926" AFTER 29480 ns,
x"00000000" AFTER 29500 ns,
x"EE6B292A" AFTER 29520 ns,
x"00000000" AFTER 29540 ns,
x"EE6B292E" AFTER 29560 ns,
x"00000000" AFTER 29580 ns,
x"EE6B2932" AFTER 29600 ns,
x"00000000" AFTER 29620 ns,
x"EE6B2936" AFTER 29640 ns,
x"00000000" AFTER 29660 ns,
x"EE6B293A" AFTER 29680 ns,
x"00000000" AFTER 29700 ns,
x"EE6B293E" AFTER 29720 ns,
x"00000000" AFTER 29740 ns,
x"EE6B2942" AFTER 29760 ns,
x"00000000" AFTER 29780 ns,
x"EE6B2946" AFTER 29800 ns,
x"00000000" AFTER 29820 ns,
x"EE6B294A" AFTER 29840 ns,
x"00000000" AFTER 29860 ns,
x"EE6B294E" AFTER 29880 ns,
x"00000000" AFTER 29900 ns,
x"EE6B2952" AFTER 29920 ns,
x"00000000" AFTER 29940 ns,
x"EE6B2956" AFTER 29960 ns,
x"00000000" AFTER 29980 ns,
x"EE6B295A" AFTER 30000 ns,
x"00000000" AFTER 30020 ns,
x"EE6B295E" AFTER 30040 ns,
x"00000000" AFTER 30060 ns,
x"EE6B2962" AFTER 30080 ns,
x"00000000" AFTER 30100 ns,
x"EE6B2966" AFTER 30120 ns,
x"00000000" AFTER 30140 ns,
x"EE6B296A" AFTER 30160 ns,
x"00000000" AFTER 30180 ns,
x"EE6B296E" AFTER 30200 ns,
x"00000000" AFTER 30220 ns,
x"EE6B2972" AFTER 30240 ns,
x"00000000" AFTER 30260 ns,
x"EE6B2976" AFTER 30280 ns,
x"00000000" AFTER 30300 ns,
x"EE6B297A" AFTER 30320 ns,
x"00000000" AFTER 30340 ns,
x"EE6B297E" AFTER 30360 ns,
x"00000000" AFTER 30380 ns,
x"EE6B2982" AFTER 30400 ns,
x"00000000" AFTER 30420 ns,
x"EE6B2986" AFTER 30440 ns,
x"00000000" AFTER 30460 ns,
x"EE6B298A" AFTER 30480 ns,
x"00000000" AFTER 30500 ns,
x"EE6B298E" AFTER 30520 ns,
x"00000000" AFTER 30540 ns,
x"EE6B2992" AFTER 30560 ns,
x"00000000" AFTER 30580 ns,
x"EE6B2996" AFTER 30600 ns,
x"00000000" AFTER 30620 ns,
x"EE6B299A" AFTER 30640 ns,
x"00000000" AFTER 30660 ns,
x"EE6B299E" AFTER 30680 ns,
x"00000000" AFTER 30700 ns,
x"EE6B29A2" AFTER 30720 ns,
x"00000000" AFTER 30740 ns,
x"EE6B29A6" AFTER 30760 ns,
x"00000000" AFTER 30780 ns,
x"EE6B29AA" AFTER 30800 ns,
x"00000000" AFTER 30820 ns,
x"EE6B29AE" AFTER 30840 ns,
x"00000000" AFTER 30860 ns,
x"EE6B29B2" AFTER 30880 ns,
x"00000000" AFTER 30900 ns,
x"EE6B29B6" AFTER 30920 ns,
x"00000000" AFTER 30940 ns,
x"EE6B29BA" AFTER 30960 ns;

PcRegisters <= x"00000000" AFTER 00020 ns,
x"00000531" AFTER 00040 ns,
x"00000000" AFTER 00060 ns,
x"0000052D" AFTER 00080 ns,
x"00000000" AFTER 00100 ns,
x"00000529" AFTER 00120 ns,
x"00000000" AFTER 00140 ns,
x"00000525" AFTER 00160 ns,
x"00000000" AFTER 00180 ns,
x"00000521" AFTER 00200 ns,
x"00000000" AFTER 00220 ns,
x"0000051D" AFTER 00240 ns,
x"00000000" AFTER 00260 ns,
x"00000519" AFTER 00280 ns,
x"00000000" AFTER 00300 ns,
x"00000515" AFTER 00320 ns,
x"00000000" AFTER 00340 ns,
x"00000511" AFTER 00360 ns,
x"00000000" AFTER 00380 ns,
x"0000050D" AFTER 00400 ns,
x"00000000" AFTER 00420 ns,
x"00000509" AFTER 00440 ns,
x"00000000" AFTER 00460 ns,
x"00000505" AFTER 00480 ns,
x"00000000" AFTER 00500 ns,
x"00000501" AFTER 00520 ns,
x"00000000" AFTER 00540 ns,
x"000004FD" AFTER 00560 ns,
x"00000000" AFTER 00580 ns,
x"000004F9" AFTER 00600 ns,
x"00000000" AFTER 00620 ns,
x"000004F5" AFTER 00640 ns,
x"00000000" AFTER 00660 ns,
x"000004F1" AFTER 00680 ns,
x"00000000" AFTER 00700 ns,
x"000004ED" AFTER 00720 ns,
x"00000000" AFTER 00740 ns,
x"000004E9" AFTER 00760 ns,
x"00000000" AFTER 00780 ns,
x"000004E5" AFTER 00800 ns,
x"00000000" AFTER 00820 ns,
x"000004E1" AFTER 00840 ns,
x"00000000" AFTER 00860 ns,
x"000004DD" AFTER 00880 ns,
x"00000000" AFTER 00900 ns,
x"000004D9" AFTER 00920 ns,
x"00000000" AFTER 00940 ns,
x"000004D5" AFTER 00960 ns,
x"00000000" AFTER 00980 ns,
x"000004D1" AFTER 01000 ns,
x"00000000" AFTER 01020 ns,
x"000004CD" AFTER 01040 ns,
x"00000000" AFTER 01060 ns,
x"000004C9" AFTER 01080 ns,
x"00000000" AFTER 01100 ns,
x"000004C5" AFTER 01120 ns,
x"00000000" AFTER 01140 ns,
x"000004C1" AFTER 01160 ns,
x"00000000" AFTER 01180 ns,
x"000004BD" AFTER 01200 ns,
x"00000000" AFTER 01220 ns,
x"000004B9" AFTER 01240 ns,
x"00000000" AFTER 01260 ns,
x"000004B5" AFTER 01280 ns,
x"00000000" AFTER 01300 ns,
x"000004B1" AFTER 01320 ns,
x"00000000" AFTER 01340 ns,
x"000004AD" AFTER 01360 ns,
x"00000000" AFTER 01380 ns,
x"000004A9" AFTER 01400 ns,
x"00000000" AFTER 01420 ns,
x"000004A5" AFTER 01440 ns,
x"00000000" AFTER 01460 ns,
x"000004A1" AFTER 01480 ns,
x"00000000" AFTER 01500 ns,
x"0000049D" AFTER 01520 ns,
x"00000000" AFTER 01540 ns,
x"00000499" AFTER 01560 ns,
x"00000000" AFTER 01580 ns,
x"00000495" AFTER 01600 ns,
x"00000000" AFTER 01620 ns,
x"00000491" AFTER 01640 ns,
x"00000000" AFTER 01660 ns,
x"0000048D" AFTER 01680 ns,
x"00000000" AFTER 01700 ns,
x"00000489" AFTER 01720 ns,
x"00000000" AFTER 01740 ns,
x"00000485" AFTER 01760 ns,
x"00000000" AFTER 01780 ns,
x"00000481" AFTER 01800 ns,
x"00000000" AFTER 01820 ns,
x"0000047D" AFTER 01840 ns,
x"00000000" AFTER 01860 ns,
x"00000479" AFTER 01880 ns,
x"00000000" AFTER 01900 ns,
x"00000475" AFTER 01920 ns,
x"00000000" AFTER 01940 ns,
x"00000471" AFTER 01960 ns,
x"00000000" AFTER 01980 ns,
x"0000046D" AFTER 02000 ns,
x"00000000" AFTER 02020 ns,
x"00000469" AFTER 02040 ns,
x"00000000" AFTER 02060 ns,
x"00000465" AFTER 02080 ns,
x"00000000" AFTER 02100 ns,
x"00000461" AFTER 02120 ns,
x"00000000" AFTER 02140 ns,
x"0000045D" AFTER 02160 ns,
x"00000000" AFTER 02180 ns,
x"00000459" AFTER 02200 ns,
x"00000000" AFTER 02220 ns,
x"00000455" AFTER 02240 ns,
x"00000000" AFTER 02260 ns,
x"00000451" AFTER 02280 ns,
x"00000000" AFTER 02300 ns,
x"0000044D" AFTER 02320 ns,
x"00000000" AFTER 02340 ns,
x"00000449" AFTER 02360 ns,
x"00000000" AFTER 02380 ns,
x"00000445" AFTER 02400 ns,
x"00000000" AFTER 02420 ns,
x"00000441" AFTER 02440 ns,
x"00000000" AFTER 02460 ns,
x"0000043D" AFTER 02480 ns,
x"00000000" AFTER 02500 ns,
x"00000439" AFTER 02520 ns,
x"00000000" AFTER 02540 ns,
x"00000435" AFTER 02560 ns,
x"00000000" AFTER 02580 ns,
x"00000431" AFTER 02600 ns,
x"00000000" AFTER 02620 ns,
x"0000042D" AFTER 02640 ns,
x"00000000" AFTER 02660 ns,
x"00000429" AFTER 02680 ns,
x"00000000" AFTER 02700 ns,
x"00000425" AFTER 02720 ns,
x"00000000" AFTER 02740 ns,
x"00000421" AFTER 02760 ns,
x"00000000" AFTER 02780 ns,
x"0000041D" AFTER 02800 ns,
x"00000000" AFTER 02820 ns,
x"00000419" AFTER 02840 ns,
x"00000000" AFTER 02860 ns,
x"00000415" AFTER 02880 ns,
x"00000000" AFTER 02900 ns,
x"00000411" AFTER 02920 ns,
x"00000000" AFTER 02940 ns,
x"0000040D" AFTER 02960 ns,
x"00000000" AFTER 02980 ns,
x"00000409" AFTER 03000 ns,
x"00000000" AFTER 03020 ns,
x"00000405" AFTER 03040 ns,
x"00000000" AFTER 03060 ns,
x"00000401" AFTER 03080 ns,
x"00000000" AFTER 03100 ns,
x"000003FD" AFTER 03120 ns,
x"00000000" AFTER 03140 ns,
x"000003F9" AFTER 03160 ns,
x"00000000" AFTER 03180 ns,
x"000003F5" AFTER 03200 ns,
x"00000000" AFTER 03220 ns,
x"000003F1" AFTER 03240 ns,
x"00000000" AFTER 03260 ns,
x"000003ED" AFTER 03280 ns,
x"00000000" AFTER 03300 ns,
x"000003E9" AFTER 03320 ns,
x"00000000" AFTER 03340 ns,
x"000003E5" AFTER 03360 ns,
x"00000000" AFTER 03380 ns,
x"000003E1" AFTER 03400 ns,
x"00000000" AFTER 03420 ns,
x"000003DD" AFTER 03440 ns,
x"00000000" AFTER 03460 ns,
x"000003D9" AFTER 03480 ns,
x"00000000" AFTER 03500 ns,
x"000003D5" AFTER 03520 ns,
x"00000000" AFTER 03540 ns,
x"000003D1" AFTER 03560 ns,
x"00000000" AFTER 03580 ns,
x"000003CD" AFTER 03600 ns,
x"00000000" AFTER 03620 ns,
x"000003C9" AFTER 03640 ns,
x"00000000" AFTER 03660 ns,
x"000003C5" AFTER 03680 ns,
x"00000000" AFTER 03700 ns,
x"000003C1" AFTER 03720 ns,
x"00000000" AFTER 03740 ns,
x"000003BD" AFTER 03760 ns,
x"00000000" AFTER 03780 ns,
x"000003B9" AFTER 03800 ns,
x"00000000" AFTER 03820 ns,
x"000003B5" AFTER 03840 ns,
x"00000000" AFTER 03860 ns,
x"000003B1" AFTER 03880 ns,
x"00000000" AFTER 03900 ns,
x"000003AD" AFTER 03920 ns,
x"00000000" AFTER 03940 ns,
x"000003A9" AFTER 03960 ns,
x"00000000" AFTER 03980 ns,
x"000003A5" AFTER 04000 ns,
x"00000000" AFTER 04020 ns,
x"000003A1" AFTER 04040 ns,
x"00000000" AFTER 04060 ns,
x"0000039D" AFTER 04080 ns,
x"00000000" AFTER 04100 ns,
x"00000399" AFTER 04120 ns,
x"00000000" AFTER 04140 ns,
x"00000395" AFTER 04160 ns,
x"00000000" AFTER 04180 ns,
x"00000391" AFTER 04200 ns,
x"00000000" AFTER 04220 ns,
x"0000038D" AFTER 04240 ns,
x"00000000" AFTER 04260 ns,
x"00000389" AFTER 04280 ns,
x"00000000" AFTER 04300 ns,
x"00000385" AFTER 04320 ns,
x"00000000" AFTER 04340 ns,
x"00000381" AFTER 04360 ns,
x"00000000" AFTER 04380 ns,
x"0000037D" AFTER 04400 ns,
x"00000000" AFTER 04420 ns,
x"00000379" AFTER 04440 ns,
x"00000000" AFTER 04460 ns,
x"00000375" AFTER 04480 ns,
x"00000000" AFTER 04500 ns,
x"00000371" AFTER 04520 ns,
x"00000000" AFTER 04540 ns,
x"0000036D" AFTER 04560 ns,
x"00000000" AFTER 04580 ns,
x"00000369" AFTER 04600 ns,
x"00000000" AFTER 04620 ns,
x"00000365" AFTER 04640 ns,
x"00000000" AFTER 04660 ns,
x"00000361" AFTER 04680 ns,
x"00000000" AFTER 04700 ns,
x"0000035D" AFTER 04720 ns,
x"00000000" AFTER 04740 ns,
x"00000359" AFTER 04760 ns,
x"00000000" AFTER 04780 ns,
x"00000355" AFTER 04800 ns,
x"00000000" AFTER 04820 ns,
x"00000351" AFTER 04840 ns,
x"00000000" AFTER 04860 ns,
x"0000034D" AFTER 04880 ns,
x"00000000" AFTER 04900 ns,
x"00000349" AFTER 04920 ns,
x"00000000" AFTER 04940 ns,
x"00000345" AFTER 04960 ns,
x"00000000" AFTER 04980 ns,
x"00000341" AFTER 05000 ns,
x"00000000" AFTER 05020 ns,
x"0000033D" AFTER 05040 ns,
x"00000000" AFTER 05060 ns,
x"00000339" AFTER 05080 ns,
x"00000000" AFTER 05100 ns,
x"00000335" AFTER 05120 ns,
x"00000000" AFTER 05140 ns,
x"00000331" AFTER 05160 ns,
x"00000000" AFTER 05180 ns,
x"0000032D" AFTER 05200 ns,
x"00000000" AFTER 05220 ns,
x"00000329" AFTER 05240 ns,
x"00000000" AFTER 05260 ns,
x"00000325" AFTER 05280 ns,
x"00000000" AFTER 05300 ns,
x"00000321" AFTER 05320 ns,
x"00000000" AFTER 05340 ns,
x"0000031D" AFTER 05360 ns,
x"00000000" AFTER 05380 ns,
x"00000319" AFTER 05400 ns,
x"00000000" AFTER 05420 ns,
x"00000315" AFTER 05440 ns,
x"00000000" AFTER 05460 ns,
x"00000311" AFTER 05480 ns,
x"00000000" AFTER 05500 ns,
x"0000030D" AFTER 05520 ns,
x"00000000" AFTER 05540 ns,
x"00000309" AFTER 05560 ns,
x"00000000" AFTER 05580 ns,
x"00000305" AFTER 05600 ns,
x"00000000" AFTER 05620 ns,
x"00000301" AFTER 05640 ns,
x"00000000" AFTER 05660 ns,
x"000002FD" AFTER 05680 ns,
x"00000000" AFTER 05700 ns,
x"000002F9" AFTER 05720 ns,
x"00000000" AFTER 05740 ns,
x"000002F5" AFTER 05760 ns,
x"00000000" AFTER 05780 ns,
x"000002F1" AFTER 05800 ns,
x"00000000" AFTER 05820 ns,
x"000002ED" AFTER 05840 ns,
x"00000000" AFTER 05860 ns,
x"000002E9" AFTER 05880 ns,
x"00000000" AFTER 05900 ns,
x"000002E5" AFTER 05920 ns,
x"00000000" AFTER 05940 ns,
x"000002E1" AFTER 05960 ns,
x"00000000" AFTER 05980 ns,
x"000002DD" AFTER 06000 ns,
x"00000000" AFTER 06020 ns,
x"000002D9" AFTER 06040 ns,
x"00000000" AFTER 06060 ns,
x"000002D5" AFTER 06080 ns,
x"00000000" AFTER 06100 ns,
x"000002D1" AFTER 06120 ns,
x"00000000" AFTER 06140 ns,
x"000002CD" AFTER 06160 ns,
x"00000000" AFTER 06180 ns,
x"000002C9" AFTER 06200 ns,
x"00000000" AFTER 06220 ns,
x"000002C5" AFTER 06240 ns,
x"00000000" AFTER 06260 ns,
x"000002C1" AFTER 06280 ns,
x"00000000" AFTER 06300 ns,
x"000002BD" AFTER 06320 ns,
x"00000000" AFTER 06340 ns,
x"000002B9" AFTER 06360 ns,
x"00000000" AFTER 06380 ns,
x"000002B5" AFTER 06400 ns,
x"00000000" AFTER 06420 ns,
x"000002B1" AFTER 06440 ns,
x"00000000" AFTER 06460 ns,
x"000002AD" AFTER 06480 ns,
x"00000000" AFTER 06500 ns,
x"000002A9" AFTER 06520 ns,
x"00000000" AFTER 06540 ns,
x"000002A5" AFTER 06560 ns,
x"00000000" AFTER 06580 ns,
x"000002A1" AFTER 06600 ns,
x"00000000" AFTER 06620 ns,
x"0000029D" AFTER 06640 ns,
x"00000000" AFTER 06660 ns,
x"00000299" AFTER 06680 ns,
x"00000000" AFTER 06700 ns,
x"00000295" AFTER 06720 ns,
x"00000000" AFTER 06740 ns,
x"00000291" AFTER 06760 ns,
x"00000000" AFTER 06780 ns,
x"0000028D" AFTER 06800 ns,
x"00000000" AFTER 06820 ns,
x"00000289" AFTER 06840 ns,
x"00000000" AFTER 06860 ns,
x"00000285" AFTER 06880 ns,
x"00000000" AFTER 06900 ns,
x"00000281" AFTER 06920 ns,
x"00000000" AFTER 06940 ns,
x"0000027D" AFTER 06960 ns,
x"00000000" AFTER 06980 ns,
x"00000279" AFTER 07000 ns,
x"00000000" AFTER 07020 ns,
x"00000275" AFTER 07040 ns,
x"00000000" AFTER 07060 ns,
x"00000271" AFTER 07080 ns,
x"00000000" AFTER 07100 ns,
x"0000026D" AFTER 07120 ns,
x"00000000" AFTER 07140 ns,
x"00000269" AFTER 07160 ns,
x"00000000" AFTER 07180 ns,
x"00000265" AFTER 07200 ns,
x"00000000" AFTER 07220 ns,
x"00000261" AFTER 07240 ns,
x"00000000" AFTER 07260 ns,
x"0000025D" AFTER 07280 ns,
x"00000000" AFTER 07300 ns,
x"00000259" AFTER 07320 ns,
x"00000000" AFTER 07340 ns,
x"00000255" AFTER 07360 ns,
x"00000000" AFTER 07380 ns,
x"00000251" AFTER 07400 ns,
x"00000000" AFTER 07420 ns,
x"0000024D" AFTER 07440 ns,
x"00000000" AFTER 07460 ns,
x"00000249" AFTER 07480 ns,
x"00000000" AFTER 07500 ns,
x"00000245" AFTER 07520 ns,
x"00000000" AFTER 07540 ns,
x"00000241" AFTER 07560 ns,
x"00000000" AFTER 07580 ns,
x"0000023D" AFTER 07600 ns,
x"00000000" AFTER 07620 ns,
x"00000239" AFTER 07640 ns,
x"00000000" AFTER 07660 ns,
x"00000235" AFTER 07680 ns,
x"00000000" AFTER 07700 ns,
x"00000231" AFTER 07720 ns,
x"00000000" AFTER 07740 ns,
x"0000022D" AFTER 07760 ns,
x"00000000" AFTER 07780 ns,
x"00000229" AFTER 07800 ns,
x"00000000" AFTER 07820 ns,
x"00000225" AFTER 07840 ns,
x"00000000" AFTER 07860 ns,
x"00000221" AFTER 07880 ns,
x"00000000" AFTER 07900 ns,
x"0000021D" AFTER 07920 ns,
x"00000000" AFTER 07940 ns,
x"00000219" AFTER 07960 ns,
x"00000000" AFTER 07980 ns,
x"00000215" AFTER 08000 ns,
x"00000000" AFTER 08020 ns,
x"00000211" AFTER 08040 ns,
x"00000000" AFTER 08060 ns,
x"0000020D" AFTER 08080 ns,
x"00000000" AFTER 08100 ns,
x"00000209" AFTER 08120 ns,
x"00000000" AFTER 08140 ns,
x"00000205" AFTER 08160 ns,
x"00000000" AFTER 08180 ns,
x"00000201" AFTER 08200 ns,
x"00000000" AFTER 08220 ns,
x"000001FD" AFTER 08240 ns,
x"00000000" AFTER 08260 ns,
x"000001F9" AFTER 08280 ns,
x"00000000" AFTER 08300 ns,
x"000001F5" AFTER 08320 ns,
x"00000000" AFTER 08340 ns,
x"000001F1" AFTER 08360 ns,
x"00000000" AFTER 08380 ns,
x"000001ED" AFTER 08400 ns,
x"00000000" AFTER 08420 ns,
x"000001E9" AFTER 08440 ns,
x"00000000" AFTER 08460 ns,
x"000001E5" AFTER 08480 ns,
x"00000000" AFTER 08500 ns,
x"000001E1" AFTER 08520 ns,
x"00000000" AFTER 08540 ns,
x"000001DD" AFTER 08560 ns,
x"00000000" AFTER 08580 ns,
x"000001D9" AFTER 08600 ns,
x"00000000" AFTER 08620 ns,
x"000001D5" AFTER 08640 ns,
x"00000000" AFTER 08660 ns,
x"000001D1" AFTER 08680 ns,
x"00000000" AFTER 08700 ns,
x"000001CD" AFTER 08720 ns,
x"00000000" AFTER 08740 ns,
x"000001C9" AFTER 08760 ns,
x"00000000" AFTER 08780 ns,
x"000001C5" AFTER 08800 ns,
x"00000000" AFTER 08820 ns,
x"000001C1" AFTER 08840 ns,
x"00000000" AFTER 08860 ns,
x"000001BD" AFTER 08880 ns,
x"00000000" AFTER 08900 ns,
x"000001B9" AFTER 08920 ns,
x"00000000" AFTER 08940 ns,
x"000001B5" AFTER 08960 ns,
x"00000000" AFTER 08980 ns,
x"000001B1" AFTER 09000 ns,
x"00000000" AFTER 09020 ns,
x"000001AD" AFTER 09040 ns,
x"00000000" AFTER 09060 ns,
x"000001A9" AFTER 09080 ns,
x"00000000" AFTER 09100 ns,
x"000001A5" AFTER 09120 ns,
x"00000000" AFTER 09140 ns,
x"000001A1" AFTER 09160 ns,
x"00000000" AFTER 09180 ns,
x"0000019D" AFTER 09200 ns,
x"00000000" AFTER 09220 ns,
x"00000199" AFTER 09240 ns,
x"00000000" AFTER 09260 ns,
x"00000195" AFTER 09280 ns,
x"00000000" AFTER 09300 ns,
x"00000191" AFTER 09320 ns,
x"00000000" AFTER 09340 ns,
x"0000018D" AFTER 09360 ns,
x"00000000" AFTER 09380 ns,
x"00000189" AFTER 09400 ns,
x"00000000" AFTER 09420 ns,
x"00000185" AFTER 09440 ns,
x"00000000" AFTER 09460 ns,
x"00000181" AFTER 09480 ns,
x"00000000" AFTER 09500 ns,
x"0000017D" AFTER 09520 ns,
x"00000000" AFTER 09540 ns,
x"00000179" AFTER 09560 ns,
x"00000000" AFTER 09580 ns,
x"00000175" AFTER 09600 ns,
x"00000000" AFTER 09620 ns,
x"00000171" AFTER 09640 ns,
x"00000000" AFTER 09660 ns,
x"0000016D" AFTER 09680 ns,
x"00000000" AFTER 09700 ns,
x"00000169" AFTER 09720 ns,
x"00000000" AFTER 09740 ns,
x"00000165" AFTER 09760 ns,
x"00000000" AFTER 09780 ns,
x"00000161" AFTER 09800 ns,
x"00000000" AFTER 09820 ns,
x"0000015D" AFTER 09840 ns,
x"00000000" AFTER 09860 ns,
x"00000159" AFTER 09880 ns,
x"00000000" AFTER 09900 ns,
x"00000155" AFTER 09920 ns,
x"00000000" AFTER 09940 ns,
x"00000151" AFTER 09960 ns,
x"00000000" AFTER 09980 ns,
x"0000014D" AFTER 10000 ns,
x"00000000" AFTER 10020 ns,
x"00000149" AFTER 10040 ns,
x"00000000" AFTER 10060 ns,
x"00000145" AFTER 10080 ns,
x"00000000" AFTER 10100 ns,
x"00000141" AFTER 10120 ns,
x"00000000" AFTER 10140 ns,
x"0000013D" AFTER 10160 ns,
x"00000000" AFTER 10180 ns,
x"00000139" AFTER 10200 ns,
x"00000000" AFTER 10220 ns,
x"00000135" AFTER 10240 ns,
x"00000000" AFTER 10260 ns,
x"00000131" AFTER 10280 ns,
x"00000000" AFTER 10300 ns,
x"0000012D" AFTER 10320 ns,
x"00000000" AFTER 10340 ns,
x"00000129" AFTER 10360 ns,
x"00000000" AFTER 10380 ns,
x"00000125" AFTER 10400 ns,
x"00000000" AFTER 10420 ns,
x"00000121" AFTER 10440 ns,
x"00000000" AFTER 10460 ns,
x"0000011D" AFTER 10480 ns,
x"00000000" AFTER 10500 ns,
x"00000119" AFTER 10520 ns,
x"00000000" AFTER 10540 ns,
x"00000115" AFTER 10560 ns,
x"00000000" AFTER 10580 ns,
x"00000111" AFTER 10600 ns,
x"00000000" AFTER 10620 ns,
x"0000010D" AFTER 10640 ns,
x"00000000" AFTER 10660 ns,
x"00000109" AFTER 10680 ns,
x"00000000" AFTER 10700 ns,
x"00000105" AFTER 10720 ns,
x"00000000" AFTER 10740 ns,
x"00000101" AFTER 10760 ns,
x"00000000" AFTER 10780 ns,
x"000000FD" AFTER 10800 ns,
x"00000000" AFTER 10820 ns,
x"000000F9" AFTER 10840 ns,
x"00000000" AFTER 10860 ns,
x"000000F5" AFTER 10880 ns,
x"00000000" AFTER 10900 ns,
x"000000F1" AFTER 10920 ns,
x"00000000" AFTER 10940 ns,
x"000000ED" AFTER 10960 ns,
x"00000000" AFTER 10980 ns,
x"000000E9" AFTER 11000 ns,
x"00000000" AFTER 11020 ns,
x"000000E5" AFTER 11040 ns,
x"00000000" AFTER 11060 ns,
x"000000E1" AFTER 11080 ns,
x"00000000" AFTER 11100 ns,
x"000000DD" AFTER 11120 ns,
x"00000000" AFTER 11140 ns,
x"000000D9" AFTER 11160 ns,
x"00000000" AFTER 11180 ns,
x"000000D5" AFTER 11200 ns,
x"00000000" AFTER 11220 ns,
x"000000D1" AFTER 11240 ns,
x"00000000" AFTER 11260 ns,
x"000000CD" AFTER 11280 ns,
x"00000000" AFTER 11300 ns,
x"000000C9" AFTER 11320 ns,
x"00000000" AFTER 11340 ns,
x"000000C5" AFTER 11360 ns,
x"00000000" AFTER 11380 ns,
x"000000C1" AFTER 11400 ns,
x"00000000" AFTER 11420 ns,
x"000000BD" AFTER 11440 ns,
x"00000000" AFTER 11460 ns,
x"000000B9" AFTER 11480 ns,
x"00000000" AFTER 11500 ns,
x"000000B5" AFTER 11520 ns,
x"00000000" AFTER 11540 ns,
x"000000B1" AFTER 11560 ns,
x"00000000" AFTER 11580 ns,
x"000000AD" AFTER 11600 ns,
x"00000000" AFTER 11620 ns,
x"000000A9" AFTER 11640 ns,
x"00000000" AFTER 11660 ns,
x"000000A5" AFTER 11680 ns,
x"00000000" AFTER 11700 ns,
x"000000A1" AFTER 11720 ns,
x"00000000" AFTER 11740 ns,
x"0000009D" AFTER 11760 ns,
x"00000000" AFTER 11780 ns,
x"00000099" AFTER 11800 ns,
x"00000000" AFTER 11820 ns,
x"00000095" AFTER 11840 ns,
x"00000000" AFTER 11860 ns,
x"00000091" AFTER 11880 ns,
x"00000000" AFTER 11900 ns,
x"0000008D" AFTER 11920 ns,
x"00000000" AFTER 11940 ns,
x"00000089" AFTER 11960 ns,
x"00000000" AFTER 11980 ns,
x"00000085" AFTER 12000 ns,
x"00000000" AFTER 12020 ns,
x"00000081" AFTER 12040 ns,
x"00000000" AFTER 12060 ns,
x"0000007D" AFTER 12080 ns,
x"00000000" AFTER 12100 ns,
x"00000079" AFTER 12120 ns,
x"00000000" AFTER 12140 ns,
x"00000075" AFTER 12160 ns,
x"00000000" AFTER 12180 ns,
x"00000071" AFTER 12200 ns,
x"00000000" AFTER 12220 ns,
x"0000006D" AFTER 12240 ns,
x"00000000" AFTER 12260 ns,
x"00000069" AFTER 12280 ns,
x"00000000" AFTER 12300 ns,
x"00000065" AFTER 12320 ns,
x"00000000" AFTER 12340 ns,
x"00000061" AFTER 12360 ns,
x"00000000" AFTER 12380 ns,
x"0000005D" AFTER 12400 ns,
x"00000000" AFTER 12420 ns,
x"00000059" AFTER 12440 ns,
x"00000000" AFTER 12460 ns,
x"00000055" AFTER 12480 ns,
x"00000000" AFTER 12500 ns,
x"00000051" AFTER 12520 ns,
x"00000000" AFTER 12540 ns,
x"0000004D" AFTER 12560 ns,
x"00000000" AFTER 12580 ns,
x"00000049" AFTER 12600 ns,
x"00000000" AFTER 12620 ns,
x"00000045" AFTER 12640 ns,
x"00000000" AFTER 12660 ns,
x"00000041" AFTER 12680 ns,
x"00000000" AFTER 12700 ns,
x"0000003D" AFTER 12720 ns,
x"00000000" AFTER 12740 ns,
x"00000039" AFTER 12760 ns,
x"00000000" AFTER 12780 ns,
x"00000035" AFTER 12800 ns,
x"00000000" AFTER 12820 ns,
x"00000031" AFTER 12840 ns,
x"00000000" AFTER 12860 ns,
x"0000002D" AFTER 12880 ns,
x"00000000" AFTER 12900 ns,
x"00000029" AFTER 12920 ns,
x"00000000" AFTER 12940 ns,
x"00000025" AFTER 12960 ns,
x"00000000" AFTER 12980 ns,
x"00000021" AFTER 13000 ns,
x"00000000" AFTER 13020 ns,
x"0000001D" AFTER 13040 ns,
x"00000000" AFTER 13060 ns,
x"00000019" AFTER 13080 ns,
x"00000000" AFTER 13100 ns,
x"00000015" AFTER 13120 ns,
x"00000000" AFTER 13140 ns,
x"00000011" AFTER 13160 ns,
x"00000000" AFTER 13180 ns,
x"0000000D" AFTER 13200 ns,
x"00000000" AFTER 13220 ns,
x"00000009" AFTER 13240 ns,
x"00000000" AFTER 13260 ns,
x"00000005" AFTER 13280 ns,
x"00000000" AFTER 13300 ns,
x"00000001" AFTER 13320 ns,
x"00000000" AFTER 13340 ns,
x"EE6B27F9" AFTER 13360 ns,
x"00000000" AFTER 13380 ns,
x"EE6B27F5" AFTER 13400 ns,
x"00000000" AFTER 13420 ns,
x"EE6B27F1" AFTER 13440 ns,
x"00000000" AFTER 13460 ns,
x"EE6B27ED" AFTER 13480 ns,
x"00000000" AFTER 13500 ns,
x"EE6B27E9" AFTER 13520 ns,
x"00000000" AFTER 13540 ns,
x"EE6B27E5" AFTER 13560 ns,
x"00000000" AFTER 13580 ns,
x"EE6B27E1" AFTER 13600 ns,
x"00000000" AFTER 13620 ns,
x"EE6B27DD" AFTER 13640 ns,
x"00000000" AFTER 13660 ns,
x"EE6B27D9" AFTER 13680 ns,
x"00000000" AFTER 13700 ns,
x"EE6B27D5" AFTER 13720 ns,
x"00000000" AFTER 13740 ns,
x"EE6B27D1" AFTER 13760 ns,
x"00000000" AFTER 13780 ns,
x"EE6B27CD" AFTER 13800 ns,
x"00000000" AFTER 13820 ns,
x"EE6B27C9" AFTER 13840 ns,
x"00000000" AFTER 13860 ns,
x"EE6B27C5" AFTER 13880 ns,
x"00000000" AFTER 13900 ns,
x"EE6B27C1" AFTER 13920 ns,
x"00000000" AFTER 13940 ns,
x"EE6B27BD" AFTER 13960 ns,
x"00000000" AFTER 13980 ns,
x"EE6B27B9" AFTER 14000 ns,
x"00000000" AFTER 14020 ns,
x"EE6B27B5" AFTER 14040 ns,
x"00000000" AFTER 14060 ns,
x"EE6B27B1" AFTER 14080 ns,
x"00000000" AFTER 14100 ns,
x"EE6B27AD" AFTER 14120 ns,
x"00000000" AFTER 14140 ns,
x"EE6B27A9" AFTER 14160 ns,
x"00000000" AFTER 14180 ns,
x"EE6B27A5" AFTER 14200 ns,
x"00000000" AFTER 14220 ns,
x"EE6B27A1" AFTER 14240 ns,
x"00000000" AFTER 14260 ns,
x"EE6B279D" AFTER 14280 ns,
x"00000000" AFTER 14300 ns,
x"EE6B2799" AFTER 14320 ns,
x"00000000" AFTER 14340 ns,
x"EE6B2795" AFTER 14360 ns,
x"00000000" AFTER 14380 ns,
x"EE6B2791" AFTER 14400 ns,
x"00000000" AFTER 14420 ns,
x"EE6B278D" AFTER 14440 ns,
x"00000000" AFTER 14460 ns,
x"EE6B2789" AFTER 14480 ns,
x"00000000" AFTER 14500 ns,
x"EE6B2785" AFTER 14520 ns,
x"00000000" AFTER 14540 ns,
x"EE6B2781" AFTER 14560 ns,
x"00000000" AFTER 14580 ns,
x"EE6B277D" AFTER 14600 ns,
x"00000000" AFTER 14620 ns,
x"EE6B2779" AFTER 14640 ns,
x"00000000" AFTER 14660 ns,
x"EE6B2775" AFTER 14680 ns,
x"00000000" AFTER 14700 ns,
x"EE6B2771" AFTER 14720 ns,
x"00000000" AFTER 14740 ns,
x"EE6B276D" AFTER 14760 ns,
x"00000000" AFTER 14780 ns,
x"EE6B2769" AFTER 14800 ns,
x"00000000" AFTER 14820 ns,
x"EE6B2765" AFTER 14840 ns,
x"00000000" AFTER 14860 ns,
x"EE6B2761" AFTER 14880 ns,
x"00000000" AFTER 14900 ns,
x"EE6B275D" AFTER 14920 ns,
x"00000000" AFTER 14940 ns,
x"EE6B2759" AFTER 14960 ns,
x"00000000" AFTER 14980 ns,
x"EE6B2755" AFTER 15000 ns,
x"00000000" AFTER 15020 ns,
x"EE6B2751" AFTER 15040 ns,
x"00000000" AFTER 15060 ns,
x"EE6B274D" AFTER 15080 ns,
x"00000000" AFTER 15100 ns,
x"EE6B2749" AFTER 15120 ns,
x"00000000" AFTER 15140 ns,
x"EE6B2745" AFTER 15160 ns,
x"00000000" AFTER 15180 ns,
x"EE6B2741" AFTER 15200 ns,
x"00000000" AFTER 15220 ns,
x"EE6B273D" AFTER 15240 ns,
x"00000000" AFTER 15260 ns,
x"EE6B2739" AFTER 15280 ns,
x"00000000" AFTER 15300 ns,
x"EE6B2735" AFTER 15320 ns,
x"00000000" AFTER 15340 ns,
x"EE6B2731" AFTER 15360 ns,
x"00000000" AFTER 15380 ns,
x"EE6B272D" AFTER 15400 ns,
x"00000000" AFTER 15420 ns,
x"EE6B2729" AFTER 15440 ns,
x"00000000" AFTER 15460 ns,
x"EE6B2725" AFTER 15480 ns,
x"00000000" AFTER 15500 ns,
x"EE6B2721" AFTER 15520 ns,
x"00000000" AFTER 15540 ns,
x"EE6B271D" AFTER 15560 ns,
x"00000000" AFTER 15580 ns,
x"EE6B2719" AFTER 15600 ns,
x"00000000" AFTER 15620 ns,
x"EE6B2715" AFTER 15640 ns,
x"00000000" AFTER 15660 ns,
x"EE6B2711" AFTER 15680 ns,
x"00000000" AFTER 15700 ns,
x"EE6B270D" AFTER 15720 ns,
x"00000000" AFTER 15740 ns,
x"EE6B2709" AFTER 15760 ns,
x"00000000" AFTER 15780 ns,
x"EE6B2705" AFTER 15800 ns,
x"00000000" AFTER 15820 ns,
x"EE6B2701" AFTER 15840 ns,
x"00000000" AFTER 15860 ns,
x"EE6B26FD" AFTER 15880 ns,
x"00000000" AFTER 15900 ns,
x"EE6B26F9" AFTER 15920 ns,
x"00000000" AFTER 15940 ns,
x"EE6B26F5" AFTER 15960 ns,
x"00000000" AFTER 15980 ns,
x"EE6B26F1" AFTER 16000 ns,
x"00000000" AFTER 16020 ns,
x"EE6B26ED" AFTER 16040 ns,
x"00000000" AFTER 16060 ns,
x"EE6B26E9" AFTER 16080 ns,
x"00000000" AFTER 16100 ns,
x"EE6B26E5" AFTER 16120 ns,
x"00000000" AFTER 16140 ns,
x"EE6B26E1" AFTER 16160 ns,
x"00000000" AFTER 16180 ns,
x"EE6B26DD" AFTER 16200 ns,
x"00000000" AFTER 16220 ns,
x"EE6B26D9" AFTER 16240 ns,
x"00000000" AFTER 16260 ns,
x"EE6B26D5" AFTER 16280 ns,
x"00000000" AFTER 16300 ns,
x"EE6B26D1" AFTER 16320 ns,
x"00000000" AFTER 16340 ns,
x"EE6B26CD" AFTER 16360 ns,
x"00000000" AFTER 16380 ns,
x"EE6B26C9" AFTER 16400 ns,
x"00000000" AFTER 16420 ns,
x"EE6B26C5" AFTER 16440 ns,
x"00000000" AFTER 16460 ns,
x"EE6B26C1" AFTER 16480 ns,
x"00000000" AFTER 16500 ns,
x"EE6B26BD" AFTER 16520 ns,
x"00000000" AFTER 16540 ns,
x"EE6B26B9" AFTER 16560 ns,
x"00000000" AFTER 16580 ns,
x"EE6B26B5" AFTER 16600 ns,
x"00000000" AFTER 16620 ns,
x"EE6B26B1" AFTER 16640 ns,
x"00000000" AFTER 16660 ns,
x"EE6B26AD" AFTER 16680 ns,
x"00000000" AFTER 16700 ns,
x"EE6B26A9" AFTER 16720 ns,
x"00000000" AFTER 16740 ns,
x"EE6B26A5" AFTER 16760 ns,
x"00000000" AFTER 16780 ns,
x"EE6B26A1" AFTER 16800 ns,
x"00000000" AFTER 16820 ns,
x"EE6B269D" AFTER 16840 ns,
x"00000000" AFTER 16860 ns,
x"EE6B2699" AFTER 16880 ns,
x"00000000" AFTER 16900 ns,
x"EE6B2695" AFTER 16920 ns,
x"00000000" AFTER 16940 ns,
x"EE6B2691" AFTER 16960 ns,
x"00000000" AFTER 16980 ns,
x"EE6B268D" AFTER 17000 ns,
x"00000000" AFTER 17020 ns,
x"EE6B2689" AFTER 17040 ns,
x"00000000" AFTER 17060 ns,
x"EE6B2685" AFTER 17080 ns,
x"00000000" AFTER 17100 ns,
x"EE6B2681" AFTER 17120 ns,
x"00000000" AFTER 17140 ns,
x"EE6B267D" AFTER 17160 ns,
x"00000000" AFTER 17180 ns,
x"EE6B2679" AFTER 17200 ns,
x"00000000" AFTER 17220 ns,
x"EE6B2675" AFTER 17240 ns,
x"00000000" AFTER 17260 ns,
x"EE6B2671" AFTER 17280 ns,
x"00000000" AFTER 17300 ns,
x"EE6B266D" AFTER 17320 ns,
x"00000000" AFTER 17340 ns,
x"EE6B2669" AFTER 17360 ns,
x"00000000" AFTER 17380 ns,
x"EE6B2665" AFTER 17400 ns,
x"00000000" AFTER 17420 ns,
x"EE6B2661" AFTER 17440 ns,
x"00000000" AFTER 17460 ns,
x"EE6B265D" AFTER 17480 ns,
x"00000000" AFTER 17500 ns,
x"EE6B2659" AFTER 17520 ns,
x"00000000" AFTER 17540 ns,
x"EE6B2655" AFTER 17560 ns,
x"00000000" AFTER 17580 ns,
x"EE6B2651" AFTER 17600 ns,
x"00000000" AFTER 17620 ns,
x"EE6B264D" AFTER 17640 ns,
x"00000000" AFTER 17660 ns,
x"EE6B2649" AFTER 17680 ns,
x"00000000" AFTER 17700 ns,
x"EE6B2645" AFTER 17720 ns,
x"00000000" AFTER 17740 ns,
x"EE6B2641" AFTER 17760 ns,
x"00000000" AFTER 17780 ns,
x"EE6B263D" AFTER 17800 ns,
x"00000000" AFTER 17820 ns,
x"EE6B2639" AFTER 17840 ns,
x"00000000" AFTER 17860 ns,
x"EE6B2635" AFTER 17880 ns,
x"00000000" AFTER 17900 ns,
x"EE6B2631" AFTER 17920 ns,
x"00000000" AFTER 17940 ns,
x"EE6B262D" AFTER 17960 ns,
x"00000000" AFTER 17980 ns,
x"EE6B2629" AFTER 18000 ns,
x"00000000" AFTER 18020 ns,
x"EE6B2625" AFTER 18040 ns,
x"00000000" AFTER 18060 ns,
x"EE6B2621" AFTER 18080 ns,
x"00000000" AFTER 18100 ns,
x"EE6B261D" AFTER 18120 ns,
x"00000000" AFTER 18140 ns,
x"EE6B2619" AFTER 18160 ns,
x"00000000" AFTER 18180 ns,
x"EE6B2615" AFTER 18200 ns,
x"00000000" AFTER 18220 ns,
x"EE6B2611" AFTER 18240 ns,
x"00000000" AFTER 18260 ns,
x"EE6B260D" AFTER 18280 ns,
x"00000000" AFTER 18300 ns,
x"EE6B2609" AFTER 18320 ns,
x"00000000" AFTER 18340 ns,
x"EE6B2605" AFTER 18360 ns,
x"00000000" AFTER 18380 ns,
x"EE6B2601" AFTER 18400 ns,
x"00000000" AFTER 18420 ns,
x"EE6B25FD" AFTER 18440 ns,
x"00000000" AFTER 18460 ns,
x"EE6B25F9" AFTER 18480 ns,
x"00000000" AFTER 18500 ns,
x"EE6B25F5" AFTER 18520 ns,
x"00000000" AFTER 18540 ns,
x"EE6B25F1" AFTER 18560 ns,
x"00000000" AFTER 18580 ns,
x"EE6B25ED" AFTER 18600 ns,
x"00000000" AFTER 18620 ns,
x"EE6B25E9" AFTER 18640 ns,
x"00000000" AFTER 18660 ns,
x"EE6B25E5" AFTER 18680 ns,
x"00000000" AFTER 18700 ns,
x"EE6B25E1" AFTER 18720 ns,
x"00000000" AFTER 18740 ns,
x"EE6B25DD" AFTER 18760 ns,
x"00000000" AFTER 18780 ns,
x"EE6B25D9" AFTER 18800 ns,
x"00000000" AFTER 18820 ns,
x"EE6B25D5" AFTER 18840 ns,
x"00000000" AFTER 18860 ns,
x"EE6B25D1" AFTER 18880 ns,
x"00000000" AFTER 18900 ns,
x"EE6B25CD" AFTER 18920 ns,
x"00000000" AFTER 18940 ns,
x"EE6B25C9" AFTER 18960 ns,
x"00000000" AFTER 18980 ns,
x"EE6B25C5" AFTER 19000 ns,
x"00000000" AFTER 19020 ns,
x"EE6B25C1" AFTER 19040 ns,
x"00000000" AFTER 19060 ns,
x"EE6B25BD" AFTER 19080 ns,
x"00000000" AFTER 19100 ns,
x"EE6B25B9" AFTER 19120 ns,
x"00000000" AFTER 19140 ns,
x"EE6B25B5" AFTER 19160 ns,
x"00000000" AFTER 19180 ns,
x"EE6B25B1" AFTER 19200 ns,
x"00000000" AFTER 19220 ns,
x"EE6B25AD" AFTER 19240 ns,
x"00000000" AFTER 19260 ns,
x"EE6B25A9" AFTER 19280 ns,
x"00000000" AFTER 19300 ns,
x"EE6B25A5" AFTER 19320 ns,
x"00000000" AFTER 19340 ns,
x"EE6B25A1" AFTER 19360 ns,
x"00000000" AFTER 19380 ns,
x"EE6B259D" AFTER 19400 ns,
x"00000000" AFTER 19420 ns,
x"EE6B2599" AFTER 19440 ns,
x"00000000" AFTER 19460 ns,
x"EE6B2595" AFTER 19480 ns,
x"00000000" AFTER 19500 ns,
x"EE6B2591" AFTER 19520 ns,
x"00000000" AFTER 19540 ns,
x"EE6B258D" AFTER 19560 ns,
x"00000000" AFTER 19580 ns,
x"EE6B2589" AFTER 19600 ns,
x"00000000" AFTER 19620 ns,
x"EE6B2585" AFTER 19640 ns,
x"00000000" AFTER 19660 ns,
x"EE6B2581" AFTER 19680 ns,
x"00000000" AFTER 19700 ns,
x"EE6B257D" AFTER 19720 ns,
x"00000000" AFTER 19740 ns,
x"EE6B2579" AFTER 19760 ns,
x"00000000" AFTER 19780 ns,
x"EE6B2575" AFTER 19800 ns,
x"00000000" AFTER 19820 ns,
x"EE6B2571" AFTER 19840 ns,
x"00000000" AFTER 19860 ns,
x"EE6B256D" AFTER 19880 ns,
x"00000000" AFTER 19900 ns,
x"EE6B2569" AFTER 19920 ns,
x"00000000" AFTER 19940 ns,
x"EE6B256D" AFTER 19960 ns,
x"00000000" AFTER 19980 ns,
x"EE6B2571" AFTER 20000 ns,
x"00000000" AFTER 20020 ns,
x"EE6B2575" AFTER 20040 ns,
x"00000000" AFTER 20060 ns,
x"EE6B2579" AFTER 20080 ns,
x"00000000" AFTER 20100 ns,
x"EE6B257D" AFTER 20120 ns,
x"00000000" AFTER 20140 ns,
x"EE6B2581" AFTER 20160 ns,
x"00000000" AFTER 20180 ns,
x"EE6B2585" AFTER 20200 ns,
x"00000000" AFTER 20220 ns,
x"EE6B2589" AFTER 20240 ns,
x"00000000" AFTER 20260 ns,
x"EE6B258D" AFTER 20280 ns,
x"00000000" AFTER 20300 ns,
x"EE6B2591" AFTER 20320 ns,
x"00000000" AFTER 20340 ns,
x"EE6B2595" AFTER 20360 ns,
x"00000000" AFTER 20380 ns,
x"EE6B2599" AFTER 20400 ns,
x"00000000" AFTER 20420 ns,
x"EE6B259D" AFTER 20440 ns,
x"00000000" AFTER 20460 ns,
x"EE6B25A1" AFTER 20480 ns,
x"00000000" AFTER 20500 ns,
x"EE6B25A5" AFTER 20520 ns,
x"00000000" AFTER 20540 ns,
x"EE6B25A9" AFTER 20560 ns,
x"00000000" AFTER 20580 ns,
x"EE6B25AD" AFTER 20600 ns,
x"00000000" AFTER 20620 ns,
x"EE6B25B1" AFTER 20640 ns,
x"00000000" AFTER 20660 ns,
x"EE6B25B5" AFTER 20680 ns,
x"00000000" AFTER 20700 ns,
x"EE6B25B9" AFTER 20720 ns,
x"00000000" AFTER 20740 ns,
x"EE6B25BD" AFTER 20760 ns,
x"00000000" AFTER 20780 ns,
x"EE6B25C1" AFTER 20800 ns,
x"00000000" AFTER 20820 ns,
x"EE6B25C5" AFTER 20840 ns,
x"00000000" AFTER 20860 ns,
x"EE6B25C9" AFTER 20880 ns,
x"00000000" AFTER 20900 ns,
x"EE6B25CD" AFTER 20920 ns,
x"00000000" AFTER 20940 ns,
x"EE6B25D1" AFTER 20960 ns,
x"00000000" AFTER 20980 ns,
x"EE6B25D5" AFTER 21000 ns,
x"00000000" AFTER 21020 ns,
x"EE6B25D9" AFTER 21040 ns,
x"00000000" AFTER 21060 ns,
x"EE6B25DD" AFTER 21080 ns,
x"00000000" AFTER 21100 ns,
x"EE6B25E1" AFTER 21120 ns,
x"00000000" AFTER 21140 ns,
x"EE6B25E5" AFTER 21160 ns,
x"00000000" AFTER 21180 ns,
x"EE6B25E9" AFTER 21200 ns,
x"00000000" AFTER 21220 ns,
x"EE6B25ED" AFTER 21240 ns,
x"00000000" AFTER 21260 ns,
x"EE6B25F1" AFTER 21280 ns,
x"00000000" AFTER 21300 ns,
x"EE6B25F5" AFTER 21320 ns,
x"00000000" AFTER 21340 ns,
x"EE6B25F9" AFTER 21360 ns,
x"00000000" AFTER 21380 ns,
x"EE6B25FD" AFTER 21400 ns,
x"00000000" AFTER 21420 ns,
x"EE6B2601" AFTER 21440 ns,
x"00000000" AFTER 21460 ns,
x"EE6B2605" AFTER 21480 ns,
x"00000000" AFTER 21500 ns,
x"EE6B2609" AFTER 21520 ns,
x"00000000" AFTER 21540 ns,
x"EE6B260D" AFTER 21560 ns,
x"00000000" AFTER 21580 ns,
x"EE6B2611" AFTER 21600 ns,
x"00000000" AFTER 21620 ns,
x"EE6B2615" AFTER 21640 ns,
x"00000000" AFTER 21660 ns,
x"EE6B2619" AFTER 21680 ns,
x"00000000" AFTER 21700 ns,
x"EE6B261D" AFTER 21720 ns,
x"00000000" AFTER 21740 ns,
x"EE6B2621" AFTER 21760 ns,
x"00000000" AFTER 21780 ns,
x"EE6B2625" AFTER 21800 ns,
x"00000000" AFTER 21820 ns,
x"EE6B2629" AFTER 21840 ns,
x"00000000" AFTER 21860 ns,
x"EE6B262D" AFTER 21880 ns,
x"00000000" AFTER 21900 ns,
x"EE6B2631" AFTER 21920 ns,
x"00000000" AFTER 21940 ns,
x"EE6B2635" AFTER 21960 ns,
x"00000000" AFTER 21980 ns,
x"EE6B2639" AFTER 22000 ns,
x"00000000" AFTER 22020 ns,
x"EE6B263D" AFTER 22040 ns,
x"00000000" AFTER 22060 ns,
x"EE6B2641" AFTER 22080 ns,
x"00000000" AFTER 22100 ns,
x"EE6B2645" AFTER 22120 ns,
x"00000000" AFTER 22140 ns,
x"EE6B2649" AFTER 22160 ns,
x"00000000" AFTER 22180 ns,
x"EE6B264D" AFTER 22200 ns,
x"00000000" AFTER 22220 ns,
x"EE6B2651" AFTER 22240 ns,
x"00000000" AFTER 22260 ns,
x"EE6B2655" AFTER 22280 ns,
x"00000000" AFTER 22300 ns,
x"EE6B2659" AFTER 22320 ns,
x"00000000" AFTER 22340 ns,
x"EE6B265D" AFTER 22360 ns,
x"00000000" AFTER 22380 ns,
x"EE6B2661" AFTER 22400 ns,
x"00000000" AFTER 22420 ns,
x"EE6B2665" AFTER 22440 ns,
x"00000000" AFTER 22460 ns,
x"EE6B2669" AFTER 22480 ns,
x"00000000" AFTER 22500 ns,
x"EE6B266D" AFTER 22520 ns,
x"00000000" AFTER 22540 ns,
x"EE6B2671" AFTER 22560 ns,
x"00000000" AFTER 22580 ns,
x"EE6B2675" AFTER 22600 ns,
x"00000000" AFTER 22620 ns,
x"EE6B2679" AFTER 22640 ns,
x"00000000" AFTER 22660 ns,
x"EE6B267D" AFTER 22680 ns,
x"00000000" AFTER 22700 ns,
x"EE6B2681" AFTER 22720 ns,
x"00000000" AFTER 22740 ns,
x"EE6B2685" AFTER 22760 ns,
x"00000000" AFTER 22780 ns,
x"EE6B2689" AFTER 22800 ns,
x"00000000" AFTER 22820 ns,
x"EE6B268D" AFTER 22840 ns,
x"00000000" AFTER 22860 ns,
x"EE6B2691" AFTER 22880 ns,
x"00000000" AFTER 22900 ns,
x"EE6B2695" AFTER 22920 ns,
x"00000000" AFTER 22940 ns,
x"EE6B2699" AFTER 22960 ns,
x"00000000" AFTER 22980 ns,
x"EE6B269D" AFTER 23000 ns,
x"00000000" AFTER 23020 ns,
x"EE6B26A1" AFTER 23040 ns,
x"00000000" AFTER 23060 ns,
x"EE6B26A5" AFTER 23080 ns,
x"00000000" AFTER 23100 ns,
x"EE6B26A9" AFTER 23120 ns,
x"00000000" AFTER 23140 ns,
x"EE6B26AD" AFTER 23160 ns,
x"00000000" AFTER 23180 ns,
x"EE6B26B1" AFTER 23200 ns,
x"00000000" AFTER 23220 ns,
x"EE6B26B5" AFTER 23240 ns,
x"00000000" AFTER 23260 ns,
x"EE6B26B9" AFTER 23280 ns,
x"00000000" AFTER 23300 ns,
x"EE6B26BD" AFTER 23320 ns,
x"00000000" AFTER 23340 ns,
x"EE6B26C1" AFTER 23360 ns,
x"00000000" AFTER 23380 ns,
x"EE6B26C5" AFTER 23400 ns,
x"00000000" AFTER 23420 ns,
x"EE6B26C9" AFTER 23440 ns,
x"00000000" AFTER 23460 ns,
x"EE6B26CD" AFTER 23480 ns,
x"00000000" AFTER 23500 ns,
x"EE6B26D1" AFTER 23520 ns,
x"00000000" AFTER 23540 ns,
x"EE6B26D5" AFTER 23560 ns,
x"00000000" AFTER 23580 ns,
x"EE6B26D9" AFTER 23600 ns,
x"00000000" AFTER 23620 ns,
x"EE6B26DD" AFTER 23640 ns,
x"00000000" AFTER 23660 ns,
x"EE6B26E1" AFTER 23680 ns,
x"00000000" AFTER 23700 ns,
x"EE6B26E5" AFTER 23720 ns,
x"00000000" AFTER 23740 ns,
x"EE6B26E9" AFTER 23760 ns,
x"00000000" AFTER 23780 ns,
x"EE6B26ED" AFTER 23800 ns,
x"00000000" AFTER 23820 ns,
x"EE6B26F1" AFTER 23840 ns,
x"00000000" AFTER 23860 ns,
x"EE6B26F5" AFTER 23880 ns,
x"00000000" AFTER 23900 ns,
x"EE6B26F9" AFTER 23920 ns,
x"00000000" AFTER 23940 ns,
x"EE6B26FD" AFTER 23960 ns,
x"00000000" AFTER 23980 ns,
x"EE6B2701" AFTER 24000 ns,
x"00000000" AFTER 24020 ns,
x"EE6B2705" AFTER 24040 ns,
x"00000000" AFTER 24060 ns,
x"EE6B2709" AFTER 24080 ns,
x"00000000" AFTER 24100 ns,
x"EE6B270D" AFTER 24120 ns,
x"00000000" AFTER 24140 ns,
x"EE6B2711" AFTER 24160 ns,
x"00000000" AFTER 24180 ns,
x"EE6B2715" AFTER 24200 ns,
x"00000000" AFTER 24220 ns,
x"EE6B2719" AFTER 24240 ns,
x"00000000" AFTER 24260 ns,
x"EE6B271D" AFTER 24280 ns,
x"00000000" AFTER 24300 ns,
x"EE6B2721" AFTER 24320 ns,
x"00000000" AFTER 24340 ns,
x"EE6B2725" AFTER 24360 ns,
x"00000000" AFTER 24380 ns,
x"EE6B2729" AFTER 24400 ns,
x"00000000" AFTER 24420 ns,
x"EE6B272D" AFTER 24440 ns,
x"00000000" AFTER 24460 ns,
x"EE6B2731" AFTER 24480 ns,
x"00000000" AFTER 24500 ns,
x"EE6B2735" AFTER 24520 ns,
x"00000000" AFTER 24540 ns,
x"EE6B2739" AFTER 24560 ns,
x"00000000" AFTER 24580 ns,
x"EE6B273D" AFTER 24600 ns,
x"00000000" AFTER 24620 ns,
x"EE6B2741" AFTER 24640 ns,
x"00000000" AFTER 24660 ns,
x"EE6B2745" AFTER 24680 ns,
x"00000000" AFTER 24700 ns,
x"EE6B2749" AFTER 24720 ns,
x"00000000" AFTER 24740 ns,
x"EE6B274D" AFTER 24760 ns,
x"00000000" AFTER 24780 ns,
x"EE6B2751" AFTER 24800 ns,
x"00000000" AFTER 24820 ns,
x"EE6B2755" AFTER 24840 ns,
x"00000000" AFTER 24860 ns,
x"EE6B2759" AFTER 24880 ns,
x"00000000" AFTER 24900 ns,
x"EE6B275D" AFTER 24920 ns,
x"00000000" AFTER 24940 ns,
x"EE6B2761" AFTER 24960 ns,
x"00000000" AFTER 24980 ns,
x"EE6B2765" AFTER 25000 ns,
x"00000000" AFTER 25020 ns,
x"EE6B2769" AFTER 25040 ns,
x"00000000" AFTER 25060 ns,
x"EE6B276D" AFTER 25080 ns,
x"00000000" AFTER 25100 ns,
x"EE6B2771" AFTER 25120 ns,
x"00000000" AFTER 25140 ns,
x"EE6B2775" AFTER 25160 ns,
x"00000000" AFTER 25180 ns,
x"EE6B2779" AFTER 25200 ns,
x"00000000" AFTER 25220 ns,
x"EE6B277D" AFTER 25240 ns,
x"00000000" AFTER 25260 ns,
x"EE6B2781" AFTER 25280 ns,
x"00000000" AFTER 25300 ns,
x"EE6B2785" AFTER 25320 ns,
x"00000000" AFTER 25340 ns,
x"EE6B2789" AFTER 25360 ns,
x"00000000" AFTER 25380 ns,
x"EE6B278D" AFTER 25400 ns,
x"00000000" AFTER 25420 ns,
x"EE6B2791" AFTER 25440 ns,
x"00000000" AFTER 25460 ns,
x"EE6B2795" AFTER 25480 ns,
x"00000000" AFTER 25500 ns,
x"EE6B2799" AFTER 25520 ns,
x"00000000" AFTER 25540 ns,
x"EE6B279D" AFTER 25560 ns,
x"00000000" AFTER 25580 ns,
x"EE6B27A1" AFTER 25600 ns,
x"00000000" AFTER 25620 ns,
x"EE6B27A5" AFTER 25640 ns,
x"00000000" AFTER 25660 ns,
x"EE6B27A9" AFTER 25680 ns,
x"00000000" AFTER 25700 ns,
x"EE6B27AD" AFTER 25720 ns,
x"00000000" AFTER 25740 ns,
x"EE6B27B1" AFTER 25760 ns,
x"00000000" AFTER 25780 ns,
x"EE6B27B5" AFTER 25800 ns,
x"00000000" AFTER 25820 ns,
x"EE6B27B9" AFTER 25840 ns,
x"00000000" AFTER 25860 ns,
x"EE6B27BD" AFTER 25880 ns,
x"00000000" AFTER 25900 ns,
x"EE6B27C1" AFTER 25920 ns,
x"00000000" AFTER 25940 ns,
x"EE6B27C5" AFTER 25960 ns,
x"00000000" AFTER 25980 ns,
x"EE6B27C9" AFTER 26000 ns,
x"00000000" AFTER 26020 ns,
x"EE6B27CD" AFTER 26040 ns,
x"00000000" AFTER 26060 ns,
x"EE6B27D1" AFTER 26080 ns,
x"00000000" AFTER 26100 ns,
x"EE6B27D5" AFTER 26120 ns,
x"00000000" AFTER 26140 ns,
x"EE6B27D9" AFTER 26160 ns,
x"00000000" AFTER 26180 ns,
x"EE6B27DD" AFTER 26200 ns,
x"00000000" AFTER 26220 ns,
x"EE6B27E1" AFTER 26240 ns,
x"00000000" AFTER 26260 ns,
x"EE6B27E5" AFTER 26280 ns,
x"00000000" AFTER 26300 ns,
x"EE6B27E9" AFTER 26320 ns,
x"00000000" AFTER 26340 ns,
x"EE6B27ED" AFTER 26360 ns,
x"00000000" AFTER 26380 ns,
x"EE6B27F1" AFTER 26400 ns,
x"00000000" AFTER 26420 ns,
x"EE6B27F5" AFTER 26440 ns,
x"00000000" AFTER 26460 ns,
x"EE6B27F9" AFTER 26480 ns,
x"00000000" AFTER 26500 ns,
x"EE6B27FD" AFTER 26520 ns,
x"00000000" AFTER 26540 ns,
x"EE6B2801" AFTER 26560 ns,
x"00000000" AFTER 26580 ns,
x"EE6B2805" AFTER 26600 ns,
x"00000000" AFTER 26620 ns,
x"EE6B2809" AFTER 26640 ns,
x"00000000" AFTER 26660 ns,
x"EE6B280D" AFTER 26680 ns,
x"00000000" AFTER 26700 ns,
x"EE6B2811" AFTER 26720 ns,
x"00000000" AFTER 26740 ns,
x"EE6B2815" AFTER 26760 ns,
x"00000000" AFTER 26780 ns,
x"EE6B2819" AFTER 26800 ns,
x"00000000" AFTER 26820 ns,
x"EE6B281D" AFTER 26840 ns,
x"00000000" AFTER 26860 ns,
x"EE6B2821" AFTER 26880 ns,
x"00000000" AFTER 26900 ns,
x"EE6B2825" AFTER 26920 ns,
x"00000000" AFTER 26940 ns,
x"EE6B2829" AFTER 26960 ns,
x"00000000" AFTER 26980 ns,
x"EE6B282D" AFTER 27000 ns,
x"00000000" AFTER 27020 ns,
x"EE6B2831" AFTER 27040 ns,
x"00000000" AFTER 27060 ns,
x"EE6B2835" AFTER 27080 ns,
x"00000000" AFTER 27100 ns,
x"EE6B2839" AFTER 27120 ns,
x"00000000" AFTER 27140 ns,
x"EE6B283D" AFTER 27160 ns,
x"00000000" AFTER 27180 ns,
x"EE6B2841" AFTER 27200 ns,
x"00000000" AFTER 27220 ns,
x"EE6B2845" AFTER 27240 ns,
x"00000000" AFTER 27260 ns,
x"EE6B2849" AFTER 27280 ns,
x"00000000" AFTER 27300 ns,
x"EE6B284D" AFTER 27320 ns,
x"00000000" AFTER 27340 ns,
x"EE6B2851" AFTER 27360 ns,
x"00000000" AFTER 27380 ns,
x"EE6B2855" AFTER 27400 ns,
x"00000000" AFTER 27420 ns,
x"EE6B2859" AFTER 27440 ns,
x"00000000" AFTER 27460 ns,
x"EE6B285D" AFTER 27480 ns,
x"00000000" AFTER 27500 ns,
x"EE6B2861" AFTER 27520 ns,
x"00000000" AFTER 27540 ns,
x"EE6B2865" AFTER 27560 ns,
x"00000000" AFTER 27580 ns,
x"EE6B2869" AFTER 27600 ns,
x"00000000" AFTER 27620 ns,
x"EE6B286D" AFTER 27640 ns,
x"00000000" AFTER 27660 ns,
x"EE6B2871" AFTER 27680 ns,
x"00000000" AFTER 27700 ns,
x"EE6B2875" AFTER 27720 ns,
x"00000000" AFTER 27740 ns,
x"EE6B2879" AFTER 27760 ns,
x"00000000" AFTER 27780 ns,
x"EE6B287D" AFTER 27800 ns,
x"00000000" AFTER 27820 ns,
x"EE6B2881" AFTER 27840 ns,
x"00000000" AFTER 27860 ns,
x"EE6B2885" AFTER 27880 ns,
x"00000000" AFTER 27900 ns,
x"EE6B2889" AFTER 27920 ns,
x"00000000" AFTER 27940 ns,
x"EE6B288D" AFTER 27960 ns,
x"00000000" AFTER 27980 ns,
x"EE6B2891" AFTER 28000 ns,
x"00000000" AFTER 28020 ns,
x"EE6B2895" AFTER 28040 ns,
x"00000000" AFTER 28060 ns,
x"EE6B2899" AFTER 28080 ns,
x"00000000" AFTER 28100 ns,
x"EE6B289D" AFTER 28120 ns,
x"00000000" AFTER 28140 ns,
x"EE6B28A1" AFTER 28160 ns,
x"00000000" AFTER 28180 ns,
x"EE6B28A5" AFTER 28200 ns,
x"00000000" AFTER 28220 ns,
x"EE6B28A9" AFTER 28240 ns,
x"00000000" AFTER 28260 ns,
x"EE6B28AD" AFTER 28280 ns,
x"00000000" AFTER 28300 ns,
x"EE6B28B1" AFTER 28320 ns,
x"00000000" AFTER 28340 ns,
x"EE6B28B5" AFTER 28360 ns,
x"00000000" AFTER 28380 ns,
x"EE6B28B9" AFTER 28400 ns,
x"00000000" AFTER 28420 ns,
x"EE6B28BD" AFTER 28440 ns,
x"00000000" AFTER 28460 ns,
x"EE6B28C1" AFTER 28480 ns,
x"00000000" AFTER 28500 ns,
x"EE6B28C5" AFTER 28520 ns,
x"00000000" AFTER 28540 ns,
x"EE6B28C9" AFTER 28560 ns,
x"00000000" AFTER 28580 ns,
x"EE6B28CD" AFTER 28600 ns,
x"00000000" AFTER 28620 ns,
x"EE6B28D1" AFTER 28640 ns,
x"00000000" AFTER 28660 ns,
x"EE6B28D5" AFTER 28680 ns,
x"00000000" AFTER 28700 ns,
x"EE6B28D9" AFTER 28720 ns,
x"00000000" AFTER 28740 ns,
x"EE6B28DD" AFTER 28760 ns,
x"00000000" AFTER 28780 ns,
x"EE6B28E1" AFTER 28800 ns,
x"00000000" AFTER 28820 ns,
x"EE6B28E5" AFTER 28840 ns,
x"00000000" AFTER 28860 ns,
x"EE6B28E9" AFTER 28880 ns,
x"00000000" AFTER 28900 ns,
x"EE6B28ED" AFTER 28920 ns,
x"00000000" AFTER 28940 ns,
x"EE6B28F1" AFTER 28960 ns,
x"00000000" AFTER 28980 ns,
x"EE6B28F5" AFTER 29000 ns,
x"00000000" AFTER 29020 ns,
x"EE6B28F9" AFTER 29040 ns,
x"00000000" AFTER 29060 ns,
x"EE6B28FD" AFTER 29080 ns,
x"00000000" AFTER 29100 ns,
x"EE6B2901" AFTER 29120 ns,
x"00000000" AFTER 29140 ns,
x"EE6B2905" AFTER 29160 ns,
x"00000000" AFTER 29180 ns,
x"EE6B2909" AFTER 29200 ns,
x"00000000" AFTER 29220 ns,
x"EE6B290D" AFTER 29240 ns,
x"00000000" AFTER 29260 ns,
x"EE6B2911" AFTER 29280 ns,
x"00000000" AFTER 29300 ns,
x"EE6B2915" AFTER 29320 ns,
x"00000000" AFTER 29340 ns,
x"EE6B2919" AFTER 29360 ns,
x"00000000" AFTER 29380 ns,
x"EE6B291D" AFTER 29400 ns,
x"00000000" AFTER 29420 ns,
x"EE6B2921" AFTER 29440 ns,
x"00000000" AFTER 29460 ns,
x"EE6B2925" AFTER 29480 ns,
x"00000000" AFTER 29500 ns,
x"EE6B2929" AFTER 29520 ns,
x"00000000" AFTER 29540 ns,
x"EE6B292D" AFTER 29560 ns,
x"00000000" AFTER 29580 ns,
x"EE6B2931" AFTER 29600 ns,
x"00000000" AFTER 29620 ns,
x"EE6B2935" AFTER 29640 ns,
x"00000000" AFTER 29660 ns,
x"EE6B2939" AFTER 29680 ns,
x"00000000" AFTER 29700 ns,
x"EE6B293D" AFTER 29720 ns,
x"00000000" AFTER 29740 ns,
x"EE6B2941" AFTER 29760 ns,
x"00000000" AFTER 29780 ns,
x"EE6B2945" AFTER 29800 ns,
x"00000000" AFTER 29820 ns,
x"EE6B2949" AFTER 29840 ns,
x"00000000" AFTER 29860 ns,
x"EE6B294D" AFTER 29880 ns,
x"00000000" AFTER 29900 ns,
x"EE6B2951" AFTER 29920 ns,
x"00000000" AFTER 29940 ns,
x"EE6B2955" AFTER 29960 ns,
x"00000000" AFTER 29980 ns,
x"EE6B2959" AFTER 30000 ns,
x"00000000" AFTER 30020 ns,
x"EE6B295D" AFTER 30040 ns,
x"00000000" AFTER 30060 ns,
x"EE6B2961" AFTER 30080 ns,
x"00000000" AFTER 30100 ns,
x"EE6B2965" AFTER 30120 ns,
x"00000000" AFTER 30140 ns,
x"EE6B2969" AFTER 30160 ns,
x"00000000" AFTER 30180 ns,
x"EE6B296D" AFTER 30200 ns,
x"00000000" AFTER 30220 ns,
x"EE6B2971" AFTER 30240 ns,
x"00000000" AFTER 30260 ns,
x"EE6B2975" AFTER 30280 ns,
x"00000000" AFTER 30300 ns,
x"EE6B2979" AFTER 30320 ns,
x"00000000" AFTER 30340 ns,
x"EE6B297D" AFTER 30360 ns,
x"00000000" AFTER 30380 ns,
x"EE6B2981" AFTER 30400 ns,
x"00000000" AFTER 30420 ns,
x"EE6B2985" AFTER 30440 ns,
x"00000000" AFTER 30460 ns,
x"EE6B2989" AFTER 30480 ns,
x"00000000" AFTER 30500 ns,
x"EE6B298D" AFTER 30520 ns,
x"00000000" AFTER 30540 ns,
x"EE6B2991" AFTER 30560 ns,
x"00000000" AFTER 30580 ns,
x"EE6B2995" AFTER 30600 ns,
x"00000000" AFTER 30620 ns,
x"EE6B2999" AFTER 30640 ns,
x"00000000" AFTER 30660 ns,
x"EE6B299D" AFTER 30680 ns,
x"00000000" AFTER 30700 ns,
x"EE6B29A1" AFTER 30720 ns,
x"00000000" AFTER 30740 ns,
x"EE6B29A5" AFTER 30760 ns,
x"00000000" AFTER 30780 ns,
x"EE6B29A9" AFTER 30800 ns,
x"00000000" AFTER 30820 ns,
x"EE6B29AD" AFTER 30840 ns,
x"00000000" AFTER 30860 ns,
x"EE6B29B1" AFTER 30880 ns,
x"00000000" AFTER 30900 ns,
x"EE6B29B5" AFTER 30920 ns,
x"00000000" AFTER 30940 ns,
x"EE6B29B9" AFTER 30960 ns;

END TestProtocolRegistersArch;
