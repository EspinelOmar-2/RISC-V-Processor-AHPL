--******************************************************--
--        PONTIFICIA UNIVERSIDAD JAVERIANA              --
--                Disegno Digital                       --
--          Seccion de Tecnicas Digitales               --
-- 													              --
-- Titulo :                                             --
-- Fecha  :  	D:XX M:XX Y:20XX                         --
--******************************************************--

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
LIBRARY ALTERA;
USE ALTERA.altera_primitives_components.ALL;

--******************************************************--
-- Comentarios:
--
--
--******************************************************--

ENTITY ControlUnit IS

	PORT	 (
				IrControl         : IN  STD_LOGIC_VECTOR(12 DOWNTO 0);
				CsrControl        : IN  STD_LOGIC_VECTOR( 5 DOWNTO 0);
				IRQ               : IN  STD_LOGIC_VECTOR( 3 DOWNTO 0);
				CounterControl    : IN  STD_LOGIC;
				AluControl        : IN  STD_LOGIC_VECTOR( 3 DOWNTO 0);
				Reset             : IN  STD_LOGIC;
				Clk               : IN  STD_LOGIC;
				ControlRegisters  : OUT STD_LOGIC_VECTOR(26 DOWNTO 0);
				ControlSp         : OUT STD_LOGIC_VECTOR( 1 DOWNTO 0);
				ControlPc         : OUT STD_LOGIC_VECTOR( 2 DOWNTO 0);
				ControlAlu        : OUT STD_LOGIC_VECTOR(36 DOWNTO 0);
				ControlMar        : OUT STD_LOGIC_VECTOR( 2 DOWNTO 0);
				ControlMemoryRdWr : OUT STD_LOGIC_VECTOR( 1 DOWNTO 0);
				ControlQs         : OUT STD_LOGIC_VECTOR( 6 DOWNTO 0);
				ControlError      : OUT STD_LOGIC;
				ACK               : OUT STD_LOGIC_VECTOR( 3 DOWNTO 0);
				ControlCounter    : OUT STD_LOGIC_VECTOR( 2 DOWNTO 0);
				ControlCsr        : OUT STD_LOGIC_VECTOR(18 DOWNTO 0);
				ControlIr         : OUT STD_LOGIC
			 );

END ENTITY ControlUnit;

ARCHITECTURE ControlUnitArch OF ControlUnit IS

CONSTANT HundredZero : STD_LOGIC_VECTOR(100 DOWNTO 0) := (OTHERS => '0');

SIGNAL   D           : STD_LOGIC_VECTOR(101 DOWNTO 0);
SIGNAL   Q           : STD_LOGIC_VECTOR(101 DOWNTO 0);
SIGNAL   ToState     : STD_LOGIC_VECTOR(101 DOWNTO 0);
SIGNAL   StateEx     : STD_LOGIC_VECTOR(101 DOWNTO 0);
SIGNAL   Ir          : STD_LOGIC_VECTOR( 12 DOWNTO 0);
SIGNAL   NIr         : STD_LOGIC_VECTOR( 12 DOWNTO 0);
SIGNAL   Mul         : STD_LOGIC;
SIGNAL   NIrq        : STD_LOGIC_VECTOR(  3 DOWNTO 0);
SIGNAL   Mst04       : STD_LOGIC;
SIGNAL   Mie31       : STD_LOGIC;
SIGNAL   Mie30       : STD_LOGIC;
SIGNAL   Mie29       : STD_LOGIC;
SIGNAL   Mie28       : STD_LOGIC;
SIGNAL   Mip31       : STD_LOGIC;
SIGNAL   NMst04      : STD_LOGIC;
SIGNAL   NMie31      : STD_LOGIC;
SIGNAL   NMie30      : STD_LOGIC;
SIGNAL   NMie29      : STD_LOGIC;
SIGNAL   NMie28      : STD_LOGIC;
SIGNAL   NMip31      : STD_LOGIC;

BEGIN

--******************************************************--
--
--
--
--******************************************************--

Ir      <=     IrControl;
NIr     <= NOT IrControl;

Mst04   <=     CsrControl(5);
Mie31   <=     CsrControl(4);
Mie30   <=     CsrControl(3);
Mie29   <=     CsrControl(2);
Mie28   <=     CsrControl(1);
Mip31   <=     CsrControl(0);

NMst04  <= NOT CsrControl(5);
NMie31  <= NOT CsrControl(4);
NMie30  <= NOT CsrControl(3);
NMie29  <= NOT CsrControl(2);
NMie28  <= NOT CsrControl(1);
NMip31  <= NOT CsrControl(0);

NIrq(0) <= NOT Irq(0);
NIrq(1) <= NOT Irq(1);
NIrq(2) <= NOT Irq(2);
NIrq(3) <= NOT Irq(3);

--*******************************************************************************************************--
--
--
--
--*******************************************************************************************************--

ToState(  1) <= (Q(  0)) OR
					 (Q( 88)) OR
					 (Q( 89) AND ((NMst04) OR
									  ( Mst04 AND ((NIrq(0) AND NIrq(1) AND NIrq(2) AND NIrq(3)           ) OR
													   ( Irq(0)                                     AND NMie28) OR
													   (NIrq(0) AND  Irq(1)                         AND NMie29) OR
													   (NIrq(0) AND NIrq(1) AND  Irq(2)             AND NMie30) OR
													   (NIrq(0) AND NIrq(1) AND NIrq(2) AND  Irq(3) AND NMie31))))) OR
					 (Q( 94)) OR
					 (Q( 98)) OR
					 (Q( 99)) OR
					 (Q(100)) OR
					 (Q(101));

--*******************************************************************************************************--
--
--
--
--*******************************************************************************************************--

--                                                                                                       -- [6543210]

ToState(  6) <= NIr(6) AND NIr(5) AND  Ir(4) AND NIr(3) AND  Ir(2) AND Ir(1) AND  Ir(0)                ; -- [0010111]
ToState(  8) <= NIr(6) AND  Ir(5) AND  Ir(4) AND NIr(3) AND  Ir(2) AND Ir(1) AND  Ir(0)                ; -- [0110111]
ToState(  9) <=  Ir(6) AND  Ir(5) AND NIr(4) AND             Ir(2) AND Ir(1) AND  Ir(0)                ; -- [110C111]
ToState( 15) <=  Ir(6) AND  Ir(5) AND NIr(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(15); -- [1100011]
ToState( 19) <=  Ir(6) AND  Ir(5) AND NIr(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(19); -- [1100011]
ToState( 21) <=  Ir(6) AND  Ir(5) AND NIr(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(21); -- [1100011]
ToState( 23) <= NIr(6) AND            NIr(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0)                ; -- [0C00011]
ToState( 38) <= NIr(6) AND NIr(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(38); -- [0010011]
ToState( 40) <= NIr(6) AND NIr(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(40); -- [0010011]
ToState( 44) <= NIr(6) AND NIr(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(44); -- [0010011]
ToState( 46) <= NIr(6) AND NIr(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(46); -- [0010011]
ToState( 47) <= NIr(6) AND NIr(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(47); -- [0010011]
ToState( 48) <= NIr(6) AND NIr(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(48); -- [0010011]
ToState( 49) <= NIr(6) AND NIr(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(49); -- [0010011]
ToState( 53) <= NIr(6) AND  Ir(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(53); -- [0110011]
ToState( 55) <= NIr(6) AND  Ir(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(55); -- [0110011]
ToState( 58) <= NIr(6) AND  Ir(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(58); -- [0110011]
ToState( 60) <= NIr(6) AND  Ir(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(60); -- [0110011]
ToState( 62) <= NIr(6) AND  Ir(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(62); -- [0110011]
ToState( 64) <= NIr(6) AND  Ir(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(64); -- [0110011]
ToState( 65) <= NIr(6) AND  Ir(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(65); -- [0110011]
ToState( 66) <= NIr(6) AND  Ir(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(66); -- [0110011]
ToState( 67) <=  Ir(6) AND  Ir(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0)                ; -- [1110011]
ToState( 74) <= NIr(6) AND  Ir(5) AND  Ir(4) AND NIr(3) AND NIr(2) AND Ir(1) AND  Ir(0) AND StateEx(74); -- [0110011]
ToState( 75) <=                                                        Ir(1) AND NIr(0) AND StateEx(75); -- [XXXXX10]
ToState( 79) <=                                                        Ir(1) AND NIr(0) AND StateEx(79); -- [XXXXX10]

--               Ir(15)     Ir(14)     Ir(13)     Ir(12)      Ir(30)     Ir(25)   -- [1111][3]
--                                                                                -- [5432][0]

StateEx( 15) <=             NIr(9) AND NIr(8)                                   ; -- [X00C][X]
StateEx( 19) <=              Ir(9) AND NIr(8)                                   ; -- [X10C][X]
StateEx( 21) <=              Ir(9) AND  Ir(8)                                   ; -- [X11C][X]
StateEx( 38) <=             NIr(9) AND NIr(8) AND NIr(7)                        ; -- [X000][X]
StateEx( 40) <=             NIr(9) AND  Ir(8) AND NIr(7)                        ; -- [X010][X]
StateEx( 44) <=             NIr(9) AND  Ir(8) AND  Ir(7)                        ; -- [X011][X]
StateEx( 46) <=              Ir(9) AND NIr(8) AND NIr(7)                        ; -- [X100][X]
StateEx( 47) <=              Ir(9) AND  Ir(8) AND NIr(7)                        ; -- [X110][X]
StateEx( 48) <=              Ir(9) AND  Ir(8) AND  Ir(7)                        ; -- [X111][X]
StateEx( 49) <=                        NIr(8) AND  Ir(7)                        ; -- [XC01][C]
StateEx( 53) <=             NIr(9) AND NIr(8) AND NIr(7) AND NIr(11) AND NIr(12); -- [X000][0]
StateEx( 55) <=             NIr(9) AND NIr(8) AND NIr(7) AND  Ir(11)            ; -- [X000][1]
StateEx( 58) <=                        NIr(8) AND  Ir(7)                        ; -- [XC01][C]
StateEx( 60) <=             NIr(9) AND  Ir(8) AND NIr(7)                        ; -- [X010][X]
StateEx( 62) <=             NIr(9) AND  Ir(8) AND  Ir(7)                        ; -- [X011][X]
StateEx( 64) <=              Ir(9) AND NIr(8) AND NIr(7)                        ; -- [X100][X]
StateEx( 65) <=              Ir(9) AND  Ir(8) AND NIr(7)                        ; -- [X110][X]
StateEx( 66) <=              Ir(9) AND  Ir(8) AND  Ir(7)                        ; -- [X111][X]
StateEx( 74) <=             NIr(9) AND NIr(8) AND NIr(7)             AND  Ir(12); -- [X000][X]
StateEx( 75) <=  Ir(10) AND  Ir(9) AND NIr(8)                                   ; -- [110X][X]
StateEx( 79) <= NIr(10) AND  Ir(9) AND NIr(8)                                   ; -- [010X][X]

--*******************************************************************************************************--
--
--
--
--*******************************************************************************************************--

ToState( 84) <= '0' WHEN ((ToState( 6) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState( 8) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState( 9) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(15) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(19) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(21) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(23) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(38) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(40) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(44) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(46) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(47) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(48) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(49) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(53) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(55) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(58) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(60) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(62) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(64) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(65) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(66) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(67) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(74) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(75) = '1') AND (Q(5) = '1')) ELSE
					 '0' WHEN ((ToState(79) = '1') AND (Q(5) = '1')) ELSE
					 '1' ;

--*******************************************************************************************************--
--
--
--
--*******************************************************************************************************--

ToState( 17) <= (Q( 16) AND ((NIr(7) AND      AluControl(1))                             OR
									  (Ir (7) AND (NOT AluControl(1)))                         )) OR
					 (Q( 20) AND ((NIr(7) AND      AluControl(2)  AND (NOT AluControl(1)))    OR
									  (Ir (7) AND (NOT AluControl(2)) AND (NOT AluControl(1))) )) OR
					 (Q( 22) AND ((NIr(7) AND (NOT AluControl(1)) AND (NOT AluControl(3)))    OR
								     (Ir (7) AND (NOT AluControl(1)  AND      AluControl(3))) ));

--*******************************************************************************************************--
--
--
--
--*******************************************************************************************************--

ToState( 27) <= NIr(9) AND NIr(8) AND NIr(7);
ToState( 28) <= NIr(9) AND NIr(8) AND  Ir(7);
ToState( 29) <= NIr(9) AND  Ir(8) AND NIr(7);
ToState( 30) <=  Ir(9) AND NIr(8) AND NIr(7);
ToState( 31) <=  Ir(9) AND NIr(8) AND  Ir(7);
ToState( 32) <=  Ir(5) AND NIr(8) AND NIr(7);
ToState( 34) <=  Ir(5) AND NIr(8) AND  Ir(7);
ToState( 36) <=  Ir(5) AND  Ir(8) AND NIr(7);

--*******************************************************************************************************--
--
--
--
--*******************************************************************************************************--

ToState(42) <= (Q(41) AND   (NOT AluControl(1)) AND (NOT AluControl(2))) OR
					(Q(45) AND   (NOT AluControl(1)) AND      AluControl(2) ) OR
					(Q(61) AND   (NOT AluControl(1)) AND (NOT AluControl(2))) OR
					(Q(63) AND   (NOT AluControl(1)) AND      AluControl(2) );

ToState(43) <= (Q(41) AND (((NOT AluControl(1)) AND      AluControl(2) ) OR
									(     AluControl(1))))                        OR
					(Q(45) AND (((NOT AluControl(1)) AND (NOT AluControl(2))) OR
									(     AluControl(1))))                        OR
					(Q(61) AND (((NOT AluControl(1)) AND      AluControl(2) ) OR
									(     AluControl(1))))                        OR
					(Q(63) AND (((NOT AluControl(1)) AND (NOT AluControl(2))) OR
									(     AluControl(1))));

--*******************************************************************************************************--
--
--
--
--*******************************************************************************************************--

ToState(50) <= (Q(49) AND  NIr(11) AND NIr( 9)) OR
					(Q(50) AND (NOT CounterControl)) OR
					(Q(58) AND  NIr( 9));

ToState(51) <= (Q(49) AND  NIr(11) AND  Ir( 9)) OR
					(Q(51) AND (NOT CounterControl)) OR
					(Q(58) AND   Ir( 9) AND NIr(11));

ToState(52) <= (Q(49) AND   Ir(11))             OR
					(Q(52) AND (NOT CounterControl)) OR
					(Q(58) AND   Ir( 9) AND  Ir(11));

ToState(59) <= (Q(50) AND      CounterControl) OR
					(Q(51) AND      CounterControl) OR
					(Q(52) AND      CounterControl) ;

--*******************************************************************************************************--
--
--
--
--*******************************************************************************************************--

ToState( 68) <= NIr(9) AND NIr(8) AND  Ir(7);
ToState( 69) <= NIr(9) AND  Ir(8) AND NIr(7);
ToState( 70) <= NIr(9) AND  Ir(8) AND  Ir(7);
ToState( 71) <=  Ir(9) AND NIr(8) AND  Ir(7);
ToState( 72) <=  Ir(9) AND  Ir(8) AND NIr(7);
ToState( 73) <=  Ir(9) AND  Ir(8) AND  Ir(7);

--*******************************************************************************************************--
--
--
--
--*******************************************************************************************************--

Mul          <= (Q(  5) AND      ToState   ( 74)) OR
					 (Q( 74) AND (NOT AluControl(  0)));

--*******************************************************************************************************--
--
--
--
--*******************************************************************************************************--

ToState( 89) <= (Q(  7)) OR
					 (Q(  8)) OR
					 (Q( 12)) OR
					 (Q( 14)) OR
					 (Q( 16)  AND ((NIr(7) AND (NOT AluControl(1)))  OR
										(Ir (7) AND      AluControl(1)))) OR
					 (Q( 18)) OR
					 (Q( 20)  AND ((NIr(7) AND (NOT AluControl(2))  AND (NOT AluControl(1)))  OR
					               (Ir (7) AND      AluControl(2)   AND (NOT AluControl(1)))  OR
										(                                         AluControl(1)))) OR
					 (Q( 22)  AND ((NIr(7) AND (NOT AluControl(1))  AND      AluControl(3))   OR
									   (Ir (7) AND (NOT AluControl(1))  AND (NOT AluControl(3)))  OR
										(                AluControl(1)))) OR
					 (Q( 27)) OR
					 (Q( 28)) OR
					 (Q( 29)) OR
					 (Q( 30)) OR
					 (Q( 31)) OR
					 (Q( 33)) OR
					 (Q( 35)) OR
					 (Q( 37)) OR
					 (Q( 39)) OR
					 (Q( 42)) OR
					 (Q( 43)) OR
					 (Q( 46)) OR
					 (Q( 47)) OR
					 (Q( 48)) OR
					 (Q( 54)) OR
					 (Q( 57)) OR
					 (Q( 59)) OR
					 (Q( 64)) OR
					 (Q( 65)) OR
					 (Q( 66)) OR
					 (Q( 68)) OR
					 (Q( 69)) OR
					 (Q( 70)) OR
					 (Q( 71)) OR
					 (Q( 72)) OR
					 (Q( 73)) OR
					 (Q( 74)  AND AluControl(0)) OR
					 (Q( 78)) OR
					 (Q( 83));

--*******************************************************************************************************--
--
--
--
--*******************************************************************************************************--

ToState( 90) <=  Mst04 AND  Irq(0)                                    AND Mie28 AND  Mip31;
ToState( 91) <=  Mst04 AND NIrq(0) AND  Irq(1)                        AND Mie29 AND  Mip31;
ToState( 92) <=  Mst04 AND NIrq(0) AND NIrq(1) AND  Irq(2)            AND Mie30 AND  Mip31;
ToState( 93) <=  Mst04 AND NIrq(0) AND NIrq(1) AND NIrq(2) AND Irq(3) AND Mie31 AND  Mip31;
ToState( 94) <=             Q(90)  OR   Q(91)  OR   Q(92)  OR  Q (93);
ToState( 95) <= (Mst04 AND  Irq(0)                                    AND Mie28 AND NMip31) OR
                (Mst04 AND NIrq(0) AND  Irq(1)                        AND Mie29 AND NMip31) OR
                (Mst04 AND NIrq(0) AND NIrq(1) AND  Irq(2)            AND Mie30 AND NMip31) OR
                (Mst04 AND NIrq(0) AND NIrq(1) AND NIrq(2) AND Irq(3) AND Mie31 AND NMip31) ;

ToState( 98) <=             Irq(0)                                    AND Mie28;
ToState( 99) <=            NIrq(0) AND  Irq(1)                        AND Mie29;
ToState(100) <=            NIrq(0) AND NIrq(1) AND  Irq(2)            AND Mie30;
ToState(101) <=            NIrq(0) AND NIrq(1) AND NIrq(2) AND Irq(3) AND Mie31;

--*******************************************************************************************************--
--
--
--
--*******************************************************************************************************--

D(  0) <=    '0';
D(  1) <=            ToState(  1);
D(  2) <= Q(  1);
D(  3) <= Q(  2);
D(  4) <= Q(  3);
D(  5) <= Q(  4);
D(  6) <= Q(  5) AND ToState(  6);
D(  7) <= Q(  6);
D(  8) <= Q(  5) AND ToState(  8);
D(  9) <= Q(  5) AND ToState(  9);
D( 10) <= Q(  9);
D( 11) <= Q( 10) AND Ir (3);
D( 12) <= Q( 11);
D( 13) <= Q( 10) AND NIr(3);
D( 14) <= Q( 13);
D( 15) <= Q(  5) AND ToState( 15);
D( 16) <= Q( 15);
D( 17) <=            ToState( 17);
D( 18) <= Q( 17);
D( 19) <= Q(  5) AND ToState( 19);
D( 20) <= Q( 19);
D( 21) <= Q(  5) AND ToState( 21);
D( 22) <= Q( 21);
D( 23) <= Q(  5) AND ToState( 23);
D( 24) <= Q( 23);
D( 25) <= Q( 24) AND NIr(5);
D( 26) <= Q( 25);
D( 27) <= Q( 26) AND ToState( 27);
D( 28) <= Q( 26) AND ToState( 28);
D( 29) <= Q( 26) AND ToState( 29);
D( 30) <= Q( 26) AND ToState( 30);
D( 31) <= Q( 26) AND ToState( 31);
D( 32) <= Q( 24) AND ToState( 32);
D( 33) <= Q( 32);
D( 34) <= Q( 24) AND ToState( 34);
D( 35) <= Q( 34);
D( 36) <= Q( 24) AND ToState( 36);
D( 37) <= Q( 36);
D( 38) <= Q(  5) AND ToState( 38);
D( 39) <= Q( 38);
D( 40) <= Q(  5) AND ToState( 40);
D( 41) <= Q( 40);
D( 42) <=            ToState( 42);
D( 43) <=            ToState( 43);
D( 44) <= Q(  5) AND ToState( 44);
D( 45) <= Q( 44);
D( 46) <= Q(  5) AND ToState( 46);
D( 47) <= Q(  5) AND ToState( 47);
D( 48) <= Q(  5) AND ToState( 48);
D( 49) <= Q(  5) AND ToState( 49);
D( 50) <=            ToState( 50);
D( 51) <=            ToState( 51);
D( 52) <=            ToState( 52);
D( 53) <= Q(  5) AND ToState( 53);
D( 54) <= Q( 53);
D( 55) <= Q(  5) AND ToState( 55);
D( 56) <= Q( 55);
D( 57) <= Q( 56);
D( 58) <= Q(  5) AND ToState( 58);
D( 59) <=            ToState( 59);
D( 60) <= Q(  5) AND ToState( 60);
D( 61) <= Q( 60);
D( 62) <= Q(  5) AND ToState( 62);
D( 63) <= Q( 62);
D( 64) <= Q(  5) AND ToState( 64);
D( 65) <= Q(  5) AND ToState( 65);
D( 66) <= Q(  5) AND ToState( 66);
D( 67) <= Q(  5) AND ToState( 67);
D( 68) <= Q( 67) AND ToState( 68);
D( 69) <= Q( 67) AND ToState( 69);
D( 70) <= Q( 67) AND ToState( 70);
D( 71) <= Q( 67) AND ToState( 71);
D( 72) <= Q( 67) AND ToState( 72);
D( 73) <= Q( 67) AND ToState( 73);
D( 74) <=            Mul         ;
D( 75) <= Q(  5) AND ToState( 75);
D( 76) <= Q( 75);
D( 77) <= Q( 76);
D( 78) <= Q( 77);
D( 79) <= Q(  5) AND ToState( 79);
D( 80) <= Q( 79);
D( 81) <= Q( 80);
D( 82) <= Q( 81);
D( 83) <= Q( 82);
D( 84) <= Q(  5) AND ToState( 84);
D( 85) <= Q( 84);
D( 86) <= Q( 85);
D( 87) <= Q( 86);
D( 88) <= Q( 87);
D( 89) <=            ToState( 89);
D( 90) <= Q( 89) AND ToState( 90);
D( 91) <= Q( 89) AND ToState( 91);
D( 92) <= Q( 89) AND ToState( 92);
D( 93) <= Q( 89) AND ToState( 93);
D( 94) <=            ToState( 94);
D( 95) <= Q( 89) AND ToState( 95);
D( 96) <= Q( 95);
D( 97) <= Q( 96);
D( 98) <= Q( 97) AND ToState( 98);
D( 99) <= Q( 97) AND ToState( 99);
D(100) <= Q( 97) AND ToState(100);
D(101) <= Q( 97) AND ToState(101);

PROCESS(Clk, Reset, D)

BEGIN

	IF(Reset = '1')THEN

		Q(0)            <= '1';
		Q(101 DOWNTO 1) <= HundredZero;

	ELSIF(Rising_Edge(Clk))THEN

		Q <= D;

	END IF;

END PROCESS;

--*******************************************************************************************************--
--
-- ControlPc(0)         <= Inc(Pc)
-- ControlPc(1)         <= Pc  <= Alu
-- ControlPc(2)         <= Pc  <= CSR
--
-- ControlMar(0)        <= Mar <= Pc
-- ControlMar(1)        <= Mar <= Alu
-- ControlMar(2)        <= Mar <= Registers
--
-- ControlMemoryRdWr(0) <= Read  enable
-- ControlMemoryRdWr(1) <= Write enable
--
-- ControlSp(0)         <= Inc(SP)
-- COntrolSp(1)         <= Dec(SP)
--
-- ControlCounter(0)    <= Inc(Counter)
-- ControlCounter(1)    <= IR
-- ControlCounter(2)    <= Registers
--
--*******************************************************************************************************--

ControlPc(0)         <= Q(  5);
ControlPc(1)         <= Q( 12) OR Q( 14) OR Q( 18);
ControlPc(2)         <= Q( 88) OR Q( 98) OR Q( 99) OR Q(100) OR Q(101);

ControlMar(0)        <= Q(  1);
ControlMar(1)        <= Q( 24) OR Q( 76) OR Q( 80);
ControlMar(2)        <= Q( 85) OR Q( 95);

ControlMemoryRdWr(0) <= Q(  2) OR Q(  3) OR Q(  4) OR Q( 25) OR Q( 26) OR Q( 27) OR
							   Q( 28) OR Q( 29) OR Q( 30) OR Q( 31) OR Q( 81) OR Q( 82) OR Q( 83);

ControlMemoryRdWr(1) <= Q( 32) OR Q( 33) OR Q( 34) OR Q( 35) OR Q( 36) OR Q( 37) OR 
								Q( 77) OR Q( 78) OR Q( 86) OR Q( 87) OR Q( 96) OR Q( 97);

ControlError         <= Q( 84);

ACK(0)               <= Q( 98);
ACK(1)               <= Q( 99);
ACK(2)               <= Q(100);
ACK(3)               <= Q(101);

ControlIr            <= Q(  4);

ControlSp(0)         <= Q( 78) OR Q( 87) OR Q( 97);
ControlSp(1)         <= Q( 79);

ControlCounter(0)    <= Q( 50) OR Q( 51) OR Q( 52);
ControlCounter(1)    <= Q( 49);
ControlCounter(2)    <= Q( 58);

ControlCsr( 0)       <= Q( 67);
ControlCsr( 1)       <= Q( 68);
ControlCsr( 2)       <= Q( 69);
ControlCsr( 3)       <= Q( 70);
ControlCsr( 4)       <= Q( 71);
ControlCsr( 5)       <= Q( 72);
ControlCsr( 6)       <= Q( 73);
ControlCsr( 7)       <= Q( 84);
ControlCsr( 8)       <= Q( 88);
ControlCsr( 9)       <= Q( 90);
ControlCsr(10)       <= Q( 91);
ControlCsr(11)       <= Q( 92);
ControlCsr(12)       <= Q( 93);
ControlCsr(13)       <= Q( 94);
ControlCsr(14)       <= Q( 95);
ControlCsr(15)       <= Q( 98);
ControlCsr(16)       <= Q( 99);
ControlCsr(17)       <= Q(100);
ControlCsr(18)       <= Q(101);

ControlRegisters( 0) <= Q(  7) OR Q( 10) OR Q( 53) OR Q( 54) OR Q( 59);
ControlRegisters( 1) <= Q(  8);
ControlRegisters( 2) <= Q( 13) OR Q( 14) OR Q( 23) OR Q( 24) OR Q( 40) OR Q( 41) OR
								Q( 44) OR Q( 45) OR Q( 49) OR Q( 50) OR Q( 51) OR Q( 52);
ControlRegisters( 3) <= Q( 15) OR Q( 16);
ControlRegisters( 4) <= Q( 19) OR Q( 20) OR Q( 21) OR Q( 22) OR Q( 53) OR Q( 54) OR
								Q( 55) OR Q( 56) OR Q( 60) OR Q( 61) OR Q( 62) OR Q( 63);
ControlRegisters( 5) <= Q( 27);
ControlRegisters( 6) <= Q( 28);
ControlRegisters( 7) <= Q( 29) OR Q( 83);
ControlRegisters( 8) <= Q( 30);
ControlRegisters( 9) <= Q( 31);
ControlRegisters(10) <= Q( 32) OR Q( 33);
ControlRegisters(11) <= Q( 34) OR Q( 35);
ControlRegisters(12) <= Q( 36) OR Q( 37);
ControlRegisters(13) <= Q( 38) OR Q( 72) OR Q( 73);
ControlRegisters(14) <= Q( 39);
ControlRegisters(15) <= Q( 42);
ControlRegisters(16) <= Q( 43);
ControlRegisters(17) <= Q( 46) OR Q( 47) OR Q( 48);
ControlRegisters(18) <= Q( 57) OR Q( 64) OR Q( 65) OR Q( 66) OR Q( 74);
ControlRegisters(19) <= Q( 67);
ControlRegisters(20) <= Q( 68);
ControlRegisters(21) <= Q( 69) OR Q( 70);
ControlRegisters(22) <= Q( 75) OR Q( 76) OR Q( 79) OR Q( 80);
ControlRegisters(23) <= Q( 77) OR Q( 78);
ControlRegisters(24) <= Q( 95);
ControlRegisters(25) <= Q( 86) OR Q( 87) OR Q( 96) OR Q( 97);
ControlRegisters(26) <= Q( 58);

ControlAlu( 0)       <= Q(  6);
ControlAlu( 1)       <= Q(  7);
ControlAlu( 2)       <= Q(  9);
ControlAlu( 3)       <= Q( 10);
ControlAlu( 4)       <= Q( 11);
ControlAlu( 5)       <= Q( 12);
ControlAlu( 6)       <= Q( 13);
ControlAlu( 7)       <= Q( 14);
ControlAlu( 8)       <= Q( 15) OR Q( 16) OR Q( 19) OR Q( 20) OR Q( 21) OR Q( 22) OR Q( 60) OR Q( 61) OR Q( 62) OR Q( 63);
ControlAlu( 9)       <= Q( 17);
ControlAlu(10)       <= Q( 18);
ControlAlu(11)       <= Q( 23) OR Q( 38);
ControlAlu(12)       <= Q( 24);
ControlAlu(13)       <= Q( 39);
ControlAlu(14)       <= Q( 40) OR Q( 41) OR Q( 44) OR Q( 45);
ControlAlu(15)       <= Q( 46);
ControlAlu(16)       <= Q( 47);
ControlAlu(17)       <= Q( 48);
ControlAlu(18)       <= Q( 50);
ControlAlu(19)       <= Q( 51);
ControlAlu(20)       <= Q( 52);
ControlAlu(21)       <= Q( 53) OR Q( 54);
ControlAlu(22)       <= Q( 57);
ControlAlu(23)       <= Q( 59);
ControlAlu(24)       <= Q( 64);
ControlAlu(25)       <= Q( 65);
ControlAlu(26)       <= Q( 66);
ControlAlu(27)       <= Q( 69);
ControlAlu(28)       <= Q( 70);
ControlAlu(29)       <= Q( 72);
ControlAlu(30)       <= Q( 73);
ControlAlu(31)       <= Q( 74);
ControlAlu(32)       <= Q( 75);
ControlAlu(33)       <= Q( 76);
ControlAlu(34)       <= Q( 79);
ControlAlu(35)       <= Q( 80);
ControlAlu(36)       <= Q( 49);

WITH Q SELECT
ControlQs <= "0000000" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001",
				 "0000001" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010",
				 "0000010" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100",
				 "0000011" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000",
				 "0000100" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000",
				 "0000101" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000",
				 "0000110" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000",
				 "0000111" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000",
				 "0001000" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
				 "0001001" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000",
				 "0001010" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000",
				 "0001011" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000",
				 "0001100" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000",
				 "0001101" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000",
				 "0001110" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000",
				 "0001111" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000",
				 "0010000" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000",
				 "0010001" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000",
				 "0010010" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000",
				 "0010011" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000",
				 "0010100" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000",
				 "0010101" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000",
				 "0010110" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000",
				 "0010111" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000",
				 "0011000" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000",
				 "0011001" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000",
				 "0011010" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000",
				 "0011011" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000",
				 "0011100" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000",
				 "0011101" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000",
				 "0011110" WHEN "000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000",
				 "0011111" WHEN "000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000",
				 "0100000" WHEN "000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000",
				 "0100001" WHEN "000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000",
				 "0100010" WHEN "000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000",
				 "0100011" WHEN "000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000",
				 "0100100" WHEN "000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000",
				 "0100101" WHEN "000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000",
				 "0100110" WHEN "000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000",
				 "0100111" WHEN "000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000",
				 "0101000" WHEN "000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000",
				 "0101001" WHEN "000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000",
				 "0101010" WHEN "000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000",
				 "0101011" WHEN "000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000",
				 "0101100" WHEN "000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
				 "0101101" WHEN "000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000",
				 "0101110" WHEN "000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000",
				 "0101111" WHEN "000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000",
				 "0110000" WHEN "000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000",
				 "0110001" WHEN "000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000",
				 "0110010" WHEN "000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000",
				 "0110011" WHEN "000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000",
				 "0110100" WHEN "000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000",
				 "0110101" WHEN "000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000",
				 "0110110" WHEN "000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000",
				 "0110111" WHEN "000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000",
				 "0111000" WHEN "000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000",
				 "0111001" WHEN "000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000",
				 "0111010" WHEN "000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000",
				 "0111011" WHEN "000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000",
				 "0111100" WHEN "000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000",
				 "0111101" WHEN "000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000",
				 "0111110" WHEN "000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000",
				 "0111111" WHEN "000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000",
				 "1000000" WHEN "000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000",
				 "1000001" WHEN "000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000",
				 "1000010" WHEN "000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000",
				 "1000011" WHEN "000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000",
				 "1000100" WHEN "000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000",
				 "1000101" WHEN "000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000",
				 "1000110" WHEN "000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000",
				 "1000111" WHEN "000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000",
				 "1001000" WHEN "000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1001001" WHEN "000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1001010" WHEN "000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1001011" WHEN "000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1001100" WHEN "000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1001101" WHEN "000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1001110" WHEN "000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1001111" WHEN "000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1010000" WHEN "000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1010001" WHEN "000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1010010" WHEN "000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1010011" WHEN "000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1010100" WHEN "000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1010101" WHEN "000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1010110" WHEN "000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1010111" WHEN "000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1011000" WHEN "000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1011001" WHEN "000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1011010" WHEN "000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1011011" WHEN "000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1011100" WHEN "000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1011101" WHEN "000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1011110" WHEN "000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1011111" WHEN "000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1100000" WHEN "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1100001" WHEN "000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1100010" WHEN "000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1100011" WHEN "001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1100100" WHEN "010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1100101" WHEN "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1100110" WHEN "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
				 "1100111" WHEN OTHERS;

--******************************************************--
--
-- Summon This Block:
--
--******************************************************--
--BlockN: ENTITY WORK.ControlUnit
--PORT MAP	  (IrControl         => SLV,
--				CsrControl        => SLV,
--				IRQ               => SLV,
--				CounterControl    => SLV,
--				AluControl        => SLV,
--				Reset             => SLV,
--				Clk               => SLV,
--				ControlRegisters  => SLV,
--				ControlSp         => SLV,
--				ControlPc         => SLV,
--				ControlAlu        => SLV,
--				ControlMar        => SLV,
--				ControlMemoryRdWr => SLV,
--				ControlQs         => SLV,
--				ControlError      => SLV,
--				Ack               => SLV,
--				ControlCounter    => SLV,
--				ControlCsr        => SLV,
--				ControlIr         => SLV
--			  );
--******************************************************--

END ControlUnitArch;
