
--Definicion de las bibliotecas 
library IEEE; 
use IEEE.std_logic_1164.all;
library ALTERA;
use ALTERA.altera_primitives_components.all;



--Declaracion de entradas y salidas del bloque--
Entity MulCounter is
port(
		--Entradas
	
		reloj: in std_logic;
		reset: in std_logic;
		enable:in std_logic;
		--Salidas
		endOfCount: out	std_logic	
	  );
end Entity MulCounter;    

architecture MulCounterArch of MulCounter is
	component dffe is
	port(
		d, clk, clrn, prn, ena: IN std_logic;
		q:OUT std_logic
	);
end component dffe;


signal q: std_logic_vector(1 downto 0);
signal auxSalida: std_logic;
signal auxEnable: std_logic_vector (1 downto 0);


begin


	--flips para contar de 0 a 3
	flip1: dffe port map(NOT q(0), reloj,not reset,'1',auxEnable (0), q(0));--Declaracion de los flipflops
	flip2: dffe port map(NOT q(1), reloj,not reset,'1',auxEnable (1), q(1));

	
	--Asigna los enable 
	auxEnable (0) <= enable;
	auxEnable (1) <= q(0) and enable;

	auxSalida<= (q(0) and q(1) );
	endOfCount <= auxSalida;

--******************************************************--
-- 
-- Summon This Block:
-- 
--******************************************************--
--BlockN: ENTITY WORK.MulCounter 
--PORT MAP	  (Reloj      => SLV,
--				Reset      => SLV,
--				Enable     => SLV,
--				EndOfCount => SLV
--			  );
--******************************************************--

End MulCounterArch;